module Queue(
  input   clock,
  input   reset,
  output  io_enq_ready,
  input   io_enq_valid,
  input   io_enq_bits,
  input   io_deq_ready,
  output  io_deq_valid,
  output  io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  ram [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_en; // @[Decoupled.scala 259:95]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 264:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  assign ram_io_deq_bits_MPORT_en = 1'h1;
  assign ram_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = 1'h0;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = io_deq_ready | empty; // @[Decoupled.scala 289:16 309:{24,39}]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram[initvar] = _RAND_0[0:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  maybe_full = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Multiplier(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input         io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output        io_deq_bits,
  input  [31:0] io_op1,
  input  [31:0] io_op2,
  output [63:0] io_res,
  input         io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  pipeMidStageInfo_clock; // @[Mul.scala 150:32]
  wire  pipeMidStageInfo_reset; // @[Mul.scala 150:32]
  wire  pipeMidStageInfo_io_enq_ready; // @[Mul.scala 150:32]
  wire  pipeMidStageInfo_io_enq_valid; // @[Mul.scala 150:32]
  wire  pipeMidStageInfo_io_enq_bits; // @[Mul.scala 150:32]
  wire  pipeMidStageInfo_io_deq_ready; // @[Mul.scala 150:32]
  wire  pipeMidStageInfo_io_deq_valid; // @[Mul.scala 150:32]
  wire  pipeMidStageInfo_io_deq_bits; // @[Mul.scala 150:32]
  wire  pipeFnlStageInfo_clock; // @[Mul.scala 151:32]
  wire  pipeFnlStageInfo_reset; // @[Mul.scala 151:32]
  wire  pipeFnlStageInfo_io_enq_ready; // @[Mul.scala 151:32]
  wire  pipeFnlStageInfo_io_enq_valid; // @[Mul.scala 151:32]
  wire  pipeFnlStageInfo_io_enq_bits; // @[Mul.scala 151:32]
  wire  pipeFnlStageInfo_io_deq_ready; // @[Mul.scala 151:32]
  wire  pipeFnlStageInfo_io_deq_valid; // @[Mul.scala 151:32]
  wire  pipeFnlStageInfo_io_deq_bits; // @[Mul.scala 151:32]
  wire [32:0] oriB = {io_op2[31],io_op2}; // @[Cat.scala 31:58]
  wire [32:0] ori2B = {io_op2, 1'h0}; // @[Mul.scala 329:24]
  wire [31:0] _negB_T_1 = 32'h0 - io_op2; // @[Mul.scala 330:22]
  wire [32:0] negB = {_negB_T_1[31],_negB_T_1}; // @[Cat.scala 31:58]
  wire [32:0] neg2B = 33'h0 - ori2B; // @[Mul.scala 331:22]
  wire [2:0] booth4 = {io_op1[1],io_op1[0],1'h0}; // @[Cat.scala 31:58]
  wire  _payload_T = booth4 == 3'h0; // @[Mul.scala 341:18]
  wire  _payload_T_3 = booth4 == 3'h1; // @[Mul.scala 342:18]
  wire  _payload_T_5 = ~oriB[32]; // @[Mul.scala 178:27]
  wire [33:0] _payload_T_7 = {1'h1,_payload_T_5,oriB[31:0]}; // @[Cat.scala 31:58]
  wire  _payload_T_8 = booth4 == 3'h2; // @[Mul.scala 343:18]
  wire  _payload_T_13 = booth4 == 3'h3; // @[Mul.scala 344:18]
  wire  _payload_T_15 = ~ori2B[32]; // @[Mul.scala 178:27]
  wire [33:0] _payload_T_17 = {1'h1,_payload_T_15,ori2B[31:0]}; // @[Cat.scala 31:58]
  wire  _payload_T_18 = booth4 == 3'h4; // @[Mul.scala 345:18]
  wire  _payload_T_20 = ~neg2B[32]; // @[Mul.scala 178:27]
  wire [33:0] _payload_T_22 = {1'h1,_payload_T_20,neg2B[31:0]}; // @[Cat.scala 31:58]
  wire  _payload_T_23 = booth4 == 3'h5; // @[Mul.scala 346:18]
  wire  _payload_T_25 = ~negB[32]; // @[Mul.scala 178:27]
  wire [33:0] _payload_T_27 = {1'h1,_payload_T_25,negB[31:0]}; // @[Cat.scala 31:58]
  wire  _payload_T_28 = booth4 == 3'h6; // @[Mul.scala 347:18]
  wire  _payload_T_33 = booth4 == 3'h7; // @[Mul.scala 348:18]
  wire [33:0] _payload_T_36 = _payload_T ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_37 = _payload_T_3 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_38 = _payload_T_8 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_39 = _payload_T_13 ? _payload_T_17 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_40 = _payload_T_18 ? _payload_T_22 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_41 = _payload_T_23 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_42 = _payload_T_28 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_43 = _payload_T_33 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_44 = _payload_T_36 | _payload_T_37; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_45 = _payload_T_44 | _payload_T_38; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_46 = _payload_T_45 | _payload_T_39; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_47 = _payload_T_46 | _payload_T_40; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_48 = _payload_T_47 | _payload_T_41; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_49 = _payload_T_48 | _payload_T_42; // @[Mux.scala 27:73]
  wire [33:0] payload = _payload_T_49 | _payload_T_43; // @[Mux.scala 27:73]
  wire  tree_0_0 = payload[0]; // @[Mul.scala 384:26]
  wire  tree_1_0 = payload[1]; // @[Mul.scala 384:26]
  wire  tree_2_0 = payload[2]; // @[Mul.scala 384:26]
  wire  tree_3_0 = payload[3]; // @[Mul.scala 384:26]
  wire  tree_4_0 = payload[4]; // @[Mul.scala 384:26]
  wire  tree_5_0 = payload[5]; // @[Mul.scala 384:26]
  wire  tree_6_0 = payload[6]; // @[Mul.scala 384:26]
  wire  tree_7_0 = payload[7]; // @[Mul.scala 384:26]
  wire  tree_8_0 = payload[8]; // @[Mul.scala 384:26]
  wire  tree_9_0 = payload[9]; // @[Mul.scala 384:26]
  wire  tree_10_0 = payload[10]; // @[Mul.scala 384:26]
  wire  tree_11_0 = payload[11]; // @[Mul.scala 384:26]
  wire  tree_12_0 = payload[12]; // @[Mul.scala 384:26]
  wire  tree_13_0 = payload[13]; // @[Mul.scala 384:26]
  wire  tree_14_0 = payload[14]; // @[Mul.scala 384:26]
  wire  tree_15_0 = payload[15]; // @[Mul.scala 384:26]
  wire  tree_16_0 = payload[16]; // @[Mul.scala 384:26]
  wire  tree_17_0 = payload[17]; // @[Mul.scala 384:26]
  wire  tree_18_0 = payload[18]; // @[Mul.scala 384:26]
  wire  tree_19_0 = payload[19]; // @[Mul.scala 384:26]
  wire  tree_20_0 = payload[20]; // @[Mul.scala 384:26]
  wire  tree_21_0 = payload[21]; // @[Mul.scala 384:26]
  wire  tree_22_0 = payload[22]; // @[Mul.scala 384:26]
  wire  tree_23_0 = payload[23]; // @[Mul.scala 384:26]
  wire  tree_24_0 = payload[24]; // @[Mul.scala 384:26]
  wire  tree_25_0 = payload[25]; // @[Mul.scala 384:26]
  wire  tree_26_0 = payload[26]; // @[Mul.scala 384:26]
  wire  tree_27_0 = payload[27]; // @[Mul.scala 384:26]
  wire  tree_28_0 = payload[28]; // @[Mul.scala 384:26]
  wire  tree_29_0 = payload[29]; // @[Mul.scala 384:26]
  wire  tree_30_0 = payload[30]; // @[Mul.scala 384:26]
  wire  tree_31_0 = payload[31]; // @[Mul.scala 384:26]
  wire  tree_32_0 = payload[32]; // @[Mul.scala 384:26]
  wire  tree_33_0 = payload[33]; // @[Mul.scala 384:26]
  wire [2:0] booth4_1 = io_op1[3:1]; // @[Mul.scala 338:131]
  wire  _payload_T_51 = booth4_1 == 3'h0; // @[Mul.scala 341:18]
  wire  _payload_T_54 = booth4_1 == 3'h1; // @[Mul.scala 342:18]
  wire  _payload_T_59 = booth4_1 == 3'h2; // @[Mul.scala 343:18]
  wire  _payload_T_64 = booth4_1 == 3'h3; // @[Mul.scala 344:18]
  wire  _payload_T_69 = booth4_1 == 3'h4; // @[Mul.scala 345:18]
  wire  _payload_T_74 = booth4_1 == 3'h5; // @[Mul.scala 346:18]
  wire  _payload_T_79 = booth4_1 == 3'h6; // @[Mul.scala 347:18]
  wire  _payload_T_84 = booth4_1 == 3'h7; // @[Mul.scala 348:18]
  wire [33:0] _payload_T_87 = _payload_T_51 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_88 = _payload_T_54 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_89 = _payload_T_59 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_90 = _payload_T_64 ? _payload_T_17 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_91 = _payload_T_69 ? _payload_T_22 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_92 = _payload_T_74 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_93 = _payload_T_79 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_94 = _payload_T_84 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_95 = _payload_T_87 | _payload_T_88; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_96 = _payload_T_95 | _payload_T_89; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_97 = _payload_T_96 | _payload_T_90; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_98 = _payload_T_97 | _payload_T_91; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_99 = _payload_T_98 | _payload_T_92; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_100 = _payload_T_99 | _payload_T_93; // @[Mux.scala 27:73]
  wire [33:0] payload_1 = _payload_T_100 | _payload_T_94; // @[Mux.scala 27:73]
  wire  tree_2_0_1 = payload_1[0]; // @[Mul.scala 384:26]
  wire  tree_3_0_1 = payload_1[1]; // @[Mul.scala 384:26]
  wire  tree_4_0_1 = payload_1[2]; // @[Mul.scala 384:26]
  wire  tree_5_0_1 = payload_1[3]; // @[Mul.scala 384:26]
  wire  tree_6_0_1 = payload_1[4]; // @[Mul.scala 384:26]
  wire  tree_7_0_1 = payload_1[5]; // @[Mul.scala 384:26]
  wire  tree_8_0_1 = payload_1[6]; // @[Mul.scala 384:26]
  wire  tree_9_0_1 = payload_1[7]; // @[Mul.scala 384:26]
  wire  tree_10_0_1 = payload_1[8]; // @[Mul.scala 384:26]
  wire  tree_11_0_1 = payload_1[9]; // @[Mul.scala 384:26]
  wire  tree_12_0_1 = payload_1[10]; // @[Mul.scala 384:26]
  wire  tree_13_0_1 = payload_1[11]; // @[Mul.scala 384:26]
  wire  tree_14_0_1 = payload_1[12]; // @[Mul.scala 384:26]
  wire  tree_15_0_1 = payload_1[13]; // @[Mul.scala 384:26]
  wire  tree_16_0_1 = payload_1[14]; // @[Mul.scala 384:26]
  wire  tree_17_0_1 = payload_1[15]; // @[Mul.scala 384:26]
  wire  tree_18_0_1 = payload_1[16]; // @[Mul.scala 384:26]
  wire  tree_19_0_1 = payload_1[17]; // @[Mul.scala 384:26]
  wire  tree_20_0_1 = payload_1[18]; // @[Mul.scala 384:26]
  wire  tree_21_0_1 = payload_1[19]; // @[Mul.scala 384:26]
  wire  tree_22_0_1 = payload_1[20]; // @[Mul.scala 384:26]
  wire  tree_23_0_1 = payload_1[21]; // @[Mul.scala 384:26]
  wire  tree_24_0_1 = payload_1[22]; // @[Mul.scala 384:26]
  wire  tree_25_0_1 = payload_1[23]; // @[Mul.scala 384:26]
  wire  tree_26_0_1 = payload_1[24]; // @[Mul.scala 384:26]
  wire  tree_27_0_1 = payload_1[25]; // @[Mul.scala 384:26]
  wire  tree_28_0_1 = payload_1[26]; // @[Mul.scala 384:26]
  wire  tree_29_0_1 = payload_1[27]; // @[Mul.scala 384:26]
  wire  tree_30_0_1 = payload_1[28]; // @[Mul.scala 384:26]
  wire  tree_31_0_1 = payload_1[29]; // @[Mul.scala 384:26]
  wire  tree_32_0_1 = payload_1[30]; // @[Mul.scala 384:26]
  wire  tree_33_0_1 = payload_1[31]; // @[Mul.scala 384:26]
  wire  tree_34_0 = payload_1[32]; // @[Mul.scala 384:26]
  wire  tree_35_0 = payload_1[33]; // @[Mul.scala 384:26]
  wire [2:0] booth4_2 = io_op1[5:3]; // @[Mul.scala 338:131]
  wire  _payload_T_102 = booth4_2 == 3'h0; // @[Mul.scala 341:18]
  wire  _payload_T_105 = booth4_2 == 3'h1; // @[Mul.scala 342:18]
  wire  _payload_T_110 = booth4_2 == 3'h2; // @[Mul.scala 343:18]
  wire  _payload_T_115 = booth4_2 == 3'h3; // @[Mul.scala 344:18]
  wire  _payload_T_120 = booth4_2 == 3'h4; // @[Mul.scala 345:18]
  wire  _payload_T_125 = booth4_2 == 3'h5; // @[Mul.scala 346:18]
  wire  _payload_T_130 = booth4_2 == 3'h6; // @[Mul.scala 347:18]
  wire  _payload_T_135 = booth4_2 == 3'h7; // @[Mul.scala 348:18]
  wire [33:0] _payload_T_138 = _payload_T_102 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_139 = _payload_T_105 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_140 = _payload_T_110 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_141 = _payload_T_115 ? _payload_T_17 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_142 = _payload_T_120 ? _payload_T_22 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_143 = _payload_T_125 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_144 = _payload_T_130 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_145 = _payload_T_135 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_146 = _payload_T_138 | _payload_T_139; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_147 = _payload_T_146 | _payload_T_140; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_148 = _payload_T_147 | _payload_T_141; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_149 = _payload_T_148 | _payload_T_142; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_150 = _payload_T_149 | _payload_T_143; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_151 = _payload_T_150 | _payload_T_144; // @[Mux.scala 27:73]
  wire [33:0] payload_2 = _payload_T_151 | _payload_T_145; // @[Mux.scala 27:73]
  wire  tree_4_0_2 = payload_2[0]; // @[Mul.scala 384:26]
  wire  tree_5_0_2 = payload_2[1]; // @[Mul.scala 384:26]
  wire  tree_6_0_2 = payload_2[2]; // @[Mul.scala 384:26]
  wire  tree_7_0_2 = payload_2[3]; // @[Mul.scala 384:26]
  wire  tree_8_0_2 = payload_2[4]; // @[Mul.scala 384:26]
  wire  tree_9_0_2 = payload_2[5]; // @[Mul.scala 384:26]
  wire  tree_10_0_2 = payload_2[6]; // @[Mul.scala 384:26]
  wire  tree_11_0_2 = payload_2[7]; // @[Mul.scala 384:26]
  wire  tree_12_0_2 = payload_2[8]; // @[Mul.scala 384:26]
  wire  tree_13_0_2 = payload_2[9]; // @[Mul.scala 384:26]
  wire  tree_14_0_2 = payload_2[10]; // @[Mul.scala 384:26]
  wire  tree_15_0_2 = payload_2[11]; // @[Mul.scala 384:26]
  wire  tree_16_0_2 = payload_2[12]; // @[Mul.scala 384:26]
  wire  tree_17_0_2 = payload_2[13]; // @[Mul.scala 384:26]
  wire  tree_18_0_2 = payload_2[14]; // @[Mul.scala 384:26]
  wire  tree_19_0_2 = payload_2[15]; // @[Mul.scala 384:26]
  wire  tree_20_0_2 = payload_2[16]; // @[Mul.scala 384:26]
  wire  tree_21_0_2 = payload_2[17]; // @[Mul.scala 384:26]
  wire  tree_22_0_2 = payload_2[18]; // @[Mul.scala 384:26]
  wire  tree_23_0_2 = payload_2[19]; // @[Mul.scala 384:26]
  wire  tree_24_0_2 = payload_2[20]; // @[Mul.scala 384:26]
  wire  tree_25_0_2 = payload_2[21]; // @[Mul.scala 384:26]
  wire  tree_26_0_2 = payload_2[22]; // @[Mul.scala 384:26]
  wire  tree_27_0_2 = payload_2[23]; // @[Mul.scala 384:26]
  wire  tree_28_0_2 = payload_2[24]; // @[Mul.scala 384:26]
  wire  tree_29_0_2 = payload_2[25]; // @[Mul.scala 384:26]
  wire  tree_30_0_2 = payload_2[26]; // @[Mul.scala 384:26]
  wire  tree_31_0_2 = payload_2[27]; // @[Mul.scala 384:26]
  wire  tree_32_0_2 = payload_2[28]; // @[Mul.scala 384:26]
  wire  tree_33_0_2 = payload_2[29]; // @[Mul.scala 384:26]
  wire  tree_34_0_1 = payload_2[30]; // @[Mul.scala 384:26]
  wire  tree_35_0_1 = payload_2[31]; // @[Mul.scala 384:26]
  wire  tree_36_0 = payload_2[32]; // @[Mul.scala 384:26]
  wire  tree_37_0 = payload_2[33]; // @[Mul.scala 384:26]
  wire [2:0] booth4_3 = io_op1[7:5]; // @[Mul.scala 338:131]
  wire  _payload_T_153 = booth4_3 == 3'h0; // @[Mul.scala 341:18]
  wire  _payload_T_156 = booth4_3 == 3'h1; // @[Mul.scala 342:18]
  wire  _payload_T_161 = booth4_3 == 3'h2; // @[Mul.scala 343:18]
  wire  _payload_T_166 = booth4_3 == 3'h3; // @[Mul.scala 344:18]
  wire  _payload_T_171 = booth4_3 == 3'h4; // @[Mul.scala 345:18]
  wire  _payload_T_176 = booth4_3 == 3'h5; // @[Mul.scala 346:18]
  wire  _payload_T_181 = booth4_3 == 3'h6; // @[Mul.scala 347:18]
  wire  _payload_T_186 = booth4_3 == 3'h7; // @[Mul.scala 348:18]
  wire [33:0] _payload_T_189 = _payload_T_153 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_190 = _payload_T_156 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_191 = _payload_T_161 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_192 = _payload_T_166 ? _payload_T_17 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_193 = _payload_T_171 ? _payload_T_22 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_194 = _payload_T_176 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_195 = _payload_T_181 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_196 = _payload_T_186 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_197 = _payload_T_189 | _payload_T_190; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_198 = _payload_T_197 | _payload_T_191; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_199 = _payload_T_198 | _payload_T_192; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_200 = _payload_T_199 | _payload_T_193; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_201 = _payload_T_200 | _payload_T_194; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_202 = _payload_T_201 | _payload_T_195; // @[Mux.scala 27:73]
  wire [33:0] payload_3 = _payload_T_202 | _payload_T_196; // @[Mux.scala 27:73]
  wire  tree_6_0_3 = payload_3[0]; // @[Mul.scala 384:26]
  wire  tree_7_0_3 = payload_3[1]; // @[Mul.scala 384:26]
  wire  tree_8_0_3 = payload_3[2]; // @[Mul.scala 384:26]
  wire  tree_9_0_3 = payload_3[3]; // @[Mul.scala 384:26]
  wire  tree_10_0_3 = payload_3[4]; // @[Mul.scala 384:26]
  wire  tree_11_0_3 = payload_3[5]; // @[Mul.scala 384:26]
  wire  tree_12_0_3 = payload_3[6]; // @[Mul.scala 384:26]
  wire  tree_13_0_3 = payload_3[7]; // @[Mul.scala 384:26]
  wire  tree_14_0_3 = payload_3[8]; // @[Mul.scala 384:26]
  wire  tree_15_0_3 = payload_3[9]; // @[Mul.scala 384:26]
  wire  tree_16_0_3 = payload_3[10]; // @[Mul.scala 384:26]
  wire  tree_17_0_3 = payload_3[11]; // @[Mul.scala 384:26]
  wire  tree_18_0_3 = payload_3[12]; // @[Mul.scala 384:26]
  wire  tree_19_0_3 = payload_3[13]; // @[Mul.scala 384:26]
  wire  tree_20_0_3 = payload_3[14]; // @[Mul.scala 384:26]
  wire  tree_21_0_3 = payload_3[15]; // @[Mul.scala 384:26]
  wire  tree_22_0_3 = payload_3[16]; // @[Mul.scala 384:26]
  wire  tree_23_0_3 = payload_3[17]; // @[Mul.scala 384:26]
  wire  tree_24_0_3 = payload_3[18]; // @[Mul.scala 384:26]
  wire  tree_25_0_3 = payload_3[19]; // @[Mul.scala 384:26]
  wire  tree_26_0_3 = payload_3[20]; // @[Mul.scala 384:26]
  wire  tree_27_0_3 = payload_3[21]; // @[Mul.scala 384:26]
  wire  tree_28_0_3 = payload_3[22]; // @[Mul.scala 384:26]
  wire  tree_29_0_3 = payload_3[23]; // @[Mul.scala 384:26]
  wire  tree_30_0_3 = payload_3[24]; // @[Mul.scala 384:26]
  wire  tree_31_0_3 = payload_3[25]; // @[Mul.scala 384:26]
  wire  tree_32_0_3 = payload_3[26]; // @[Mul.scala 384:26]
  wire  tree_33_0_3 = payload_3[27]; // @[Mul.scala 384:26]
  wire  tree_34_0_2 = payload_3[28]; // @[Mul.scala 384:26]
  wire  tree_35_0_2 = payload_3[29]; // @[Mul.scala 384:26]
  wire  tree_36_0_1 = payload_3[30]; // @[Mul.scala 384:26]
  wire  tree_37_0_1 = payload_3[31]; // @[Mul.scala 384:26]
  wire  tree_38_0 = payload_3[32]; // @[Mul.scala 384:26]
  wire  tree_39_0 = payload_3[33]; // @[Mul.scala 384:26]
  wire [2:0] booth4_4 = io_op1[9:7]; // @[Mul.scala 338:131]
  wire  _payload_T_204 = booth4_4 == 3'h0; // @[Mul.scala 341:18]
  wire  _payload_T_207 = booth4_4 == 3'h1; // @[Mul.scala 342:18]
  wire  _payload_T_212 = booth4_4 == 3'h2; // @[Mul.scala 343:18]
  wire  _payload_T_217 = booth4_4 == 3'h3; // @[Mul.scala 344:18]
  wire  _payload_T_222 = booth4_4 == 3'h4; // @[Mul.scala 345:18]
  wire  _payload_T_227 = booth4_4 == 3'h5; // @[Mul.scala 346:18]
  wire  _payload_T_232 = booth4_4 == 3'h6; // @[Mul.scala 347:18]
  wire  _payload_T_237 = booth4_4 == 3'h7; // @[Mul.scala 348:18]
  wire [33:0] _payload_T_240 = _payload_T_204 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_241 = _payload_T_207 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_242 = _payload_T_212 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_243 = _payload_T_217 ? _payload_T_17 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_244 = _payload_T_222 ? _payload_T_22 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_245 = _payload_T_227 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_246 = _payload_T_232 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_247 = _payload_T_237 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_248 = _payload_T_240 | _payload_T_241; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_249 = _payload_T_248 | _payload_T_242; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_250 = _payload_T_249 | _payload_T_243; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_251 = _payload_T_250 | _payload_T_244; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_252 = _payload_T_251 | _payload_T_245; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_253 = _payload_T_252 | _payload_T_246; // @[Mux.scala 27:73]
  wire [33:0] payload_4 = _payload_T_253 | _payload_T_247; // @[Mux.scala 27:73]
  wire  tree_8_0_4 = payload_4[0]; // @[Mul.scala 384:26]
  wire  tree_9_0_4 = payload_4[1]; // @[Mul.scala 384:26]
  wire  tree_10_0_4 = payload_4[2]; // @[Mul.scala 384:26]
  wire  tree_11_0_4 = payload_4[3]; // @[Mul.scala 384:26]
  wire  tree_12_0_4 = payload_4[4]; // @[Mul.scala 384:26]
  wire  tree_13_0_4 = payload_4[5]; // @[Mul.scala 384:26]
  wire  tree_14_0_4 = payload_4[6]; // @[Mul.scala 384:26]
  wire  tree_15_0_4 = payload_4[7]; // @[Mul.scala 384:26]
  wire  tree_16_0_4 = payload_4[8]; // @[Mul.scala 384:26]
  wire  tree_17_0_4 = payload_4[9]; // @[Mul.scala 384:26]
  wire  tree_18_0_4 = payload_4[10]; // @[Mul.scala 384:26]
  wire  tree_19_0_4 = payload_4[11]; // @[Mul.scala 384:26]
  wire  tree_20_0_4 = payload_4[12]; // @[Mul.scala 384:26]
  wire  tree_21_0_4 = payload_4[13]; // @[Mul.scala 384:26]
  wire  tree_22_0_4 = payload_4[14]; // @[Mul.scala 384:26]
  wire  tree_23_0_4 = payload_4[15]; // @[Mul.scala 384:26]
  wire  tree_24_0_4 = payload_4[16]; // @[Mul.scala 384:26]
  wire  tree_25_0_4 = payload_4[17]; // @[Mul.scala 384:26]
  wire  tree_26_0_4 = payload_4[18]; // @[Mul.scala 384:26]
  wire  tree_27_0_4 = payload_4[19]; // @[Mul.scala 384:26]
  wire  tree_28_0_4 = payload_4[20]; // @[Mul.scala 384:26]
  wire  tree_29_0_4 = payload_4[21]; // @[Mul.scala 384:26]
  wire  tree_30_0_4 = payload_4[22]; // @[Mul.scala 384:26]
  wire  tree_31_0_4 = payload_4[23]; // @[Mul.scala 384:26]
  wire  tree_32_0_4 = payload_4[24]; // @[Mul.scala 384:26]
  wire  tree_33_0_4 = payload_4[25]; // @[Mul.scala 384:26]
  wire  tree_34_0_3 = payload_4[26]; // @[Mul.scala 384:26]
  wire  tree_35_0_3 = payload_4[27]; // @[Mul.scala 384:26]
  wire  tree_36_0_2 = payload_4[28]; // @[Mul.scala 384:26]
  wire  tree_37_0_2 = payload_4[29]; // @[Mul.scala 384:26]
  wire  tree_38_0_1 = payload_4[30]; // @[Mul.scala 384:26]
  wire  tree_39_0_1 = payload_4[31]; // @[Mul.scala 384:26]
  wire  tree_40_0 = payload_4[32]; // @[Mul.scala 384:26]
  wire  tree_41_0 = payload_4[33]; // @[Mul.scala 384:26]
  wire [2:0] booth4_5 = io_op1[11:9]; // @[Mul.scala 338:131]
  wire  _payload_T_255 = booth4_5 == 3'h0; // @[Mul.scala 341:18]
  wire  _payload_T_258 = booth4_5 == 3'h1; // @[Mul.scala 342:18]
  wire  _payload_T_263 = booth4_5 == 3'h2; // @[Mul.scala 343:18]
  wire  _payload_T_268 = booth4_5 == 3'h3; // @[Mul.scala 344:18]
  wire  _payload_T_273 = booth4_5 == 3'h4; // @[Mul.scala 345:18]
  wire  _payload_T_278 = booth4_5 == 3'h5; // @[Mul.scala 346:18]
  wire  _payload_T_283 = booth4_5 == 3'h6; // @[Mul.scala 347:18]
  wire  _payload_T_288 = booth4_5 == 3'h7; // @[Mul.scala 348:18]
  wire [33:0] _payload_T_291 = _payload_T_255 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_292 = _payload_T_258 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_293 = _payload_T_263 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_294 = _payload_T_268 ? _payload_T_17 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_295 = _payload_T_273 ? _payload_T_22 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_296 = _payload_T_278 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_297 = _payload_T_283 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_298 = _payload_T_288 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_299 = _payload_T_291 | _payload_T_292; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_300 = _payload_T_299 | _payload_T_293; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_301 = _payload_T_300 | _payload_T_294; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_302 = _payload_T_301 | _payload_T_295; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_303 = _payload_T_302 | _payload_T_296; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_304 = _payload_T_303 | _payload_T_297; // @[Mux.scala 27:73]
  wire [33:0] payload_5 = _payload_T_304 | _payload_T_298; // @[Mux.scala 27:73]
  wire  tree_10_0_5 = payload_5[0]; // @[Mul.scala 384:26]
  wire  tree_11_0_5 = payload_5[1]; // @[Mul.scala 384:26]
  wire  tree_12_0_5 = payload_5[2]; // @[Mul.scala 384:26]
  wire  tree_13_0_5 = payload_5[3]; // @[Mul.scala 384:26]
  wire  tree_14_0_5 = payload_5[4]; // @[Mul.scala 384:26]
  wire  tree_15_0_5 = payload_5[5]; // @[Mul.scala 384:26]
  wire  tree_16_0_5 = payload_5[6]; // @[Mul.scala 384:26]
  wire  tree_17_0_5 = payload_5[7]; // @[Mul.scala 384:26]
  wire  tree_18_0_5 = payload_5[8]; // @[Mul.scala 384:26]
  wire  tree_19_0_5 = payload_5[9]; // @[Mul.scala 384:26]
  wire  tree_20_0_5 = payload_5[10]; // @[Mul.scala 384:26]
  wire  tree_21_0_5 = payload_5[11]; // @[Mul.scala 384:26]
  wire  tree_22_0_5 = payload_5[12]; // @[Mul.scala 384:26]
  wire  tree_23_0_5 = payload_5[13]; // @[Mul.scala 384:26]
  wire  tree_24_0_5 = payload_5[14]; // @[Mul.scala 384:26]
  wire  tree_25_0_5 = payload_5[15]; // @[Mul.scala 384:26]
  wire  tree_26_0_5 = payload_5[16]; // @[Mul.scala 384:26]
  wire  tree_27_0_5 = payload_5[17]; // @[Mul.scala 384:26]
  wire  tree_28_0_5 = payload_5[18]; // @[Mul.scala 384:26]
  wire  tree_29_0_5 = payload_5[19]; // @[Mul.scala 384:26]
  wire  tree_30_0_5 = payload_5[20]; // @[Mul.scala 384:26]
  wire  tree_31_0_5 = payload_5[21]; // @[Mul.scala 384:26]
  wire  tree_32_0_5 = payload_5[22]; // @[Mul.scala 384:26]
  wire  tree_33_0_5 = payload_5[23]; // @[Mul.scala 384:26]
  wire  tree_34_0_4 = payload_5[24]; // @[Mul.scala 384:26]
  wire  tree_35_0_4 = payload_5[25]; // @[Mul.scala 384:26]
  wire  tree_36_0_3 = payload_5[26]; // @[Mul.scala 384:26]
  wire  tree_37_0_3 = payload_5[27]; // @[Mul.scala 384:26]
  wire  tree_38_0_2 = payload_5[28]; // @[Mul.scala 384:26]
  wire  tree_39_0_2 = payload_5[29]; // @[Mul.scala 384:26]
  wire  tree_40_0_1 = payload_5[30]; // @[Mul.scala 384:26]
  wire  tree_41_0_1 = payload_5[31]; // @[Mul.scala 384:26]
  wire  tree_42_0 = payload_5[32]; // @[Mul.scala 384:26]
  wire  tree_43_0 = payload_5[33]; // @[Mul.scala 384:26]
  wire [2:0] booth4_6 = io_op1[13:11]; // @[Mul.scala 338:131]
  wire  _payload_T_306 = booth4_6 == 3'h0; // @[Mul.scala 341:18]
  wire  _payload_T_309 = booth4_6 == 3'h1; // @[Mul.scala 342:18]
  wire  _payload_T_314 = booth4_6 == 3'h2; // @[Mul.scala 343:18]
  wire  _payload_T_319 = booth4_6 == 3'h3; // @[Mul.scala 344:18]
  wire  _payload_T_324 = booth4_6 == 3'h4; // @[Mul.scala 345:18]
  wire  _payload_T_329 = booth4_6 == 3'h5; // @[Mul.scala 346:18]
  wire  _payload_T_334 = booth4_6 == 3'h6; // @[Mul.scala 347:18]
  wire  _payload_T_339 = booth4_6 == 3'h7; // @[Mul.scala 348:18]
  wire [33:0] _payload_T_342 = _payload_T_306 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_343 = _payload_T_309 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_344 = _payload_T_314 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_345 = _payload_T_319 ? _payload_T_17 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_346 = _payload_T_324 ? _payload_T_22 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_347 = _payload_T_329 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_348 = _payload_T_334 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_349 = _payload_T_339 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_350 = _payload_T_342 | _payload_T_343; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_351 = _payload_T_350 | _payload_T_344; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_352 = _payload_T_351 | _payload_T_345; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_353 = _payload_T_352 | _payload_T_346; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_354 = _payload_T_353 | _payload_T_347; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_355 = _payload_T_354 | _payload_T_348; // @[Mux.scala 27:73]
  wire [33:0] payload_6 = _payload_T_355 | _payload_T_349; // @[Mux.scala 27:73]
  wire  tree_12_0_6 = payload_6[0]; // @[Mul.scala 384:26]
  wire  tree_13_0_6 = payload_6[1]; // @[Mul.scala 384:26]
  wire  tree_14_0_6 = payload_6[2]; // @[Mul.scala 384:26]
  wire  tree_15_0_6 = payload_6[3]; // @[Mul.scala 384:26]
  wire  tree_16_0_6 = payload_6[4]; // @[Mul.scala 384:26]
  wire  tree_17_0_6 = payload_6[5]; // @[Mul.scala 384:26]
  wire  tree_18_0_6 = payload_6[6]; // @[Mul.scala 384:26]
  wire  tree_19_0_6 = payload_6[7]; // @[Mul.scala 384:26]
  wire  tree_20_0_6 = payload_6[8]; // @[Mul.scala 384:26]
  wire  tree_21_0_6 = payload_6[9]; // @[Mul.scala 384:26]
  wire  tree_22_0_6 = payload_6[10]; // @[Mul.scala 384:26]
  wire  tree_23_0_6 = payload_6[11]; // @[Mul.scala 384:26]
  wire  tree_24_0_6 = payload_6[12]; // @[Mul.scala 384:26]
  wire  tree_25_0_6 = payload_6[13]; // @[Mul.scala 384:26]
  wire  tree_26_0_6 = payload_6[14]; // @[Mul.scala 384:26]
  wire  tree_27_0_6 = payload_6[15]; // @[Mul.scala 384:26]
  wire  tree_28_0_6 = payload_6[16]; // @[Mul.scala 384:26]
  wire  tree_29_0_6 = payload_6[17]; // @[Mul.scala 384:26]
  wire  tree_30_0_6 = payload_6[18]; // @[Mul.scala 384:26]
  wire  tree_31_0_6 = payload_6[19]; // @[Mul.scala 384:26]
  wire  tree_32_0_6 = payload_6[20]; // @[Mul.scala 384:26]
  wire  tree_33_0_6 = payload_6[21]; // @[Mul.scala 384:26]
  wire  tree_34_0_5 = payload_6[22]; // @[Mul.scala 384:26]
  wire  tree_35_0_5 = payload_6[23]; // @[Mul.scala 384:26]
  wire  tree_36_0_4 = payload_6[24]; // @[Mul.scala 384:26]
  wire  tree_37_0_4 = payload_6[25]; // @[Mul.scala 384:26]
  wire  tree_38_0_3 = payload_6[26]; // @[Mul.scala 384:26]
  wire  tree_39_0_3 = payload_6[27]; // @[Mul.scala 384:26]
  wire  tree_40_0_2 = payload_6[28]; // @[Mul.scala 384:26]
  wire  tree_41_0_2 = payload_6[29]; // @[Mul.scala 384:26]
  wire  tree_42_0_1 = payload_6[30]; // @[Mul.scala 384:26]
  wire  tree_43_0_1 = payload_6[31]; // @[Mul.scala 384:26]
  wire  tree_44_0 = payload_6[32]; // @[Mul.scala 384:26]
  wire  tree_45_0 = payload_6[33]; // @[Mul.scala 384:26]
  wire [2:0] booth4_7 = io_op1[15:13]; // @[Mul.scala 338:131]
  wire  _payload_T_357 = booth4_7 == 3'h0; // @[Mul.scala 341:18]
  wire  _payload_T_360 = booth4_7 == 3'h1; // @[Mul.scala 342:18]
  wire  _payload_T_365 = booth4_7 == 3'h2; // @[Mul.scala 343:18]
  wire  _payload_T_370 = booth4_7 == 3'h3; // @[Mul.scala 344:18]
  wire  _payload_T_375 = booth4_7 == 3'h4; // @[Mul.scala 345:18]
  wire  _payload_T_380 = booth4_7 == 3'h5; // @[Mul.scala 346:18]
  wire  _payload_T_385 = booth4_7 == 3'h6; // @[Mul.scala 347:18]
  wire  _payload_T_390 = booth4_7 == 3'h7; // @[Mul.scala 348:18]
  wire [33:0] _payload_T_393 = _payload_T_357 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_394 = _payload_T_360 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_395 = _payload_T_365 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_396 = _payload_T_370 ? _payload_T_17 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_397 = _payload_T_375 ? _payload_T_22 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_398 = _payload_T_380 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_399 = _payload_T_385 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_400 = _payload_T_390 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_401 = _payload_T_393 | _payload_T_394; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_402 = _payload_T_401 | _payload_T_395; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_403 = _payload_T_402 | _payload_T_396; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_404 = _payload_T_403 | _payload_T_397; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_405 = _payload_T_404 | _payload_T_398; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_406 = _payload_T_405 | _payload_T_399; // @[Mux.scala 27:73]
  wire [33:0] payload_7 = _payload_T_406 | _payload_T_400; // @[Mux.scala 27:73]
  wire  tree_14_0_7 = payload_7[0]; // @[Mul.scala 384:26]
  wire  tree_15_0_7 = payload_7[1]; // @[Mul.scala 384:26]
  wire  tree_16_0_7 = payload_7[2]; // @[Mul.scala 384:26]
  wire  tree_17_0_7 = payload_7[3]; // @[Mul.scala 384:26]
  wire  tree_18_0_7 = payload_7[4]; // @[Mul.scala 384:26]
  wire  tree_19_0_7 = payload_7[5]; // @[Mul.scala 384:26]
  wire  tree_20_0_7 = payload_7[6]; // @[Mul.scala 384:26]
  wire  tree_21_0_7 = payload_7[7]; // @[Mul.scala 384:26]
  wire  tree_22_0_7 = payload_7[8]; // @[Mul.scala 384:26]
  wire  tree_23_0_7 = payload_7[9]; // @[Mul.scala 384:26]
  wire  tree_24_0_7 = payload_7[10]; // @[Mul.scala 384:26]
  wire  tree_25_0_7 = payload_7[11]; // @[Mul.scala 384:26]
  wire  tree_26_0_7 = payload_7[12]; // @[Mul.scala 384:26]
  wire  tree_27_0_7 = payload_7[13]; // @[Mul.scala 384:26]
  wire  tree_28_0_7 = payload_7[14]; // @[Mul.scala 384:26]
  wire  tree_29_0_7 = payload_7[15]; // @[Mul.scala 384:26]
  wire  tree_30_0_7 = payload_7[16]; // @[Mul.scala 384:26]
  wire  tree_31_0_7 = payload_7[17]; // @[Mul.scala 384:26]
  wire  tree_32_0_7 = payload_7[18]; // @[Mul.scala 384:26]
  wire  tree_33_0_7 = payload_7[19]; // @[Mul.scala 384:26]
  wire  tree_34_0_6 = payload_7[20]; // @[Mul.scala 384:26]
  wire  tree_35_0_6 = payload_7[21]; // @[Mul.scala 384:26]
  wire  tree_36_0_5 = payload_7[22]; // @[Mul.scala 384:26]
  wire  tree_37_0_5 = payload_7[23]; // @[Mul.scala 384:26]
  wire  tree_38_0_4 = payload_7[24]; // @[Mul.scala 384:26]
  wire  tree_39_0_4 = payload_7[25]; // @[Mul.scala 384:26]
  wire  tree_40_0_3 = payload_7[26]; // @[Mul.scala 384:26]
  wire  tree_41_0_3 = payload_7[27]; // @[Mul.scala 384:26]
  wire  tree_42_0_2 = payload_7[28]; // @[Mul.scala 384:26]
  wire  tree_43_0_2 = payload_7[29]; // @[Mul.scala 384:26]
  wire  tree_44_0_1 = payload_7[30]; // @[Mul.scala 384:26]
  wire  tree_45_0_1 = payload_7[31]; // @[Mul.scala 384:26]
  wire  tree_46_0 = payload_7[32]; // @[Mul.scala 384:26]
  wire  tree_47_0 = payload_7[33]; // @[Mul.scala 384:26]
  wire [2:0] booth4_8 = io_op1[17:15]; // @[Mul.scala 338:131]
  wire  _payload_T_408 = booth4_8 == 3'h0; // @[Mul.scala 341:18]
  wire  _payload_T_411 = booth4_8 == 3'h1; // @[Mul.scala 342:18]
  wire  _payload_T_416 = booth4_8 == 3'h2; // @[Mul.scala 343:18]
  wire  _payload_T_421 = booth4_8 == 3'h3; // @[Mul.scala 344:18]
  wire  _payload_T_426 = booth4_8 == 3'h4; // @[Mul.scala 345:18]
  wire  _payload_T_431 = booth4_8 == 3'h5; // @[Mul.scala 346:18]
  wire  _payload_T_436 = booth4_8 == 3'h6; // @[Mul.scala 347:18]
  wire  _payload_T_441 = booth4_8 == 3'h7; // @[Mul.scala 348:18]
  wire [33:0] _payload_T_444 = _payload_T_408 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_445 = _payload_T_411 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_446 = _payload_T_416 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_447 = _payload_T_421 ? _payload_T_17 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_448 = _payload_T_426 ? _payload_T_22 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_449 = _payload_T_431 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_450 = _payload_T_436 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_451 = _payload_T_441 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_452 = _payload_T_444 | _payload_T_445; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_453 = _payload_T_452 | _payload_T_446; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_454 = _payload_T_453 | _payload_T_447; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_455 = _payload_T_454 | _payload_T_448; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_456 = _payload_T_455 | _payload_T_449; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_457 = _payload_T_456 | _payload_T_450; // @[Mux.scala 27:73]
  wire [33:0] payload_8 = _payload_T_457 | _payload_T_451; // @[Mux.scala 27:73]
  wire  tree_16_0_8 = payload_8[0]; // @[Mul.scala 384:26]
  wire  tree_17_0_8 = payload_8[1]; // @[Mul.scala 384:26]
  wire  tree_18_0_8 = payload_8[2]; // @[Mul.scala 384:26]
  wire  tree_19_0_8 = payload_8[3]; // @[Mul.scala 384:26]
  wire  tree_20_0_8 = payload_8[4]; // @[Mul.scala 384:26]
  wire  tree_21_0_8 = payload_8[5]; // @[Mul.scala 384:26]
  wire  tree_22_0_8 = payload_8[6]; // @[Mul.scala 384:26]
  wire  tree_23_0_8 = payload_8[7]; // @[Mul.scala 384:26]
  wire  tree_24_0_8 = payload_8[8]; // @[Mul.scala 384:26]
  wire  tree_25_0_8 = payload_8[9]; // @[Mul.scala 384:26]
  wire  tree_26_0_8 = payload_8[10]; // @[Mul.scala 384:26]
  wire  tree_27_0_8 = payload_8[11]; // @[Mul.scala 384:26]
  wire  tree_28_0_8 = payload_8[12]; // @[Mul.scala 384:26]
  wire  tree_29_0_8 = payload_8[13]; // @[Mul.scala 384:26]
  wire  tree_30_0_8 = payload_8[14]; // @[Mul.scala 384:26]
  wire  tree_31_0_8 = payload_8[15]; // @[Mul.scala 384:26]
  wire  tree_32_0_8 = payload_8[16]; // @[Mul.scala 384:26]
  wire  tree_33_0_8 = payload_8[17]; // @[Mul.scala 384:26]
  wire  tree_34_0_7 = payload_8[18]; // @[Mul.scala 384:26]
  wire  tree_35_0_7 = payload_8[19]; // @[Mul.scala 384:26]
  wire  tree_36_0_6 = payload_8[20]; // @[Mul.scala 384:26]
  wire  tree_37_0_6 = payload_8[21]; // @[Mul.scala 384:26]
  wire  tree_38_0_5 = payload_8[22]; // @[Mul.scala 384:26]
  wire  tree_39_0_5 = payload_8[23]; // @[Mul.scala 384:26]
  wire  tree_40_0_4 = payload_8[24]; // @[Mul.scala 384:26]
  wire  tree_41_0_4 = payload_8[25]; // @[Mul.scala 384:26]
  wire  tree_42_0_3 = payload_8[26]; // @[Mul.scala 384:26]
  wire  tree_43_0_3 = payload_8[27]; // @[Mul.scala 384:26]
  wire  tree_44_0_2 = payload_8[28]; // @[Mul.scala 384:26]
  wire  tree_45_0_2 = payload_8[29]; // @[Mul.scala 384:26]
  wire  tree_46_0_1 = payload_8[30]; // @[Mul.scala 384:26]
  wire  tree_47_0_1 = payload_8[31]; // @[Mul.scala 384:26]
  wire  tree_48_0 = payload_8[32]; // @[Mul.scala 384:26]
  wire  tree_49_0 = payload_8[33]; // @[Mul.scala 384:26]
  wire [2:0] booth4_9 = io_op1[19:17]; // @[Mul.scala 338:131]
  wire  _payload_T_459 = booth4_9 == 3'h0; // @[Mul.scala 341:18]
  wire  _payload_T_462 = booth4_9 == 3'h1; // @[Mul.scala 342:18]
  wire  _payload_T_467 = booth4_9 == 3'h2; // @[Mul.scala 343:18]
  wire  _payload_T_472 = booth4_9 == 3'h3; // @[Mul.scala 344:18]
  wire  _payload_T_477 = booth4_9 == 3'h4; // @[Mul.scala 345:18]
  wire  _payload_T_482 = booth4_9 == 3'h5; // @[Mul.scala 346:18]
  wire  _payload_T_487 = booth4_9 == 3'h6; // @[Mul.scala 347:18]
  wire  _payload_T_492 = booth4_9 == 3'h7; // @[Mul.scala 348:18]
  wire [33:0] _payload_T_495 = _payload_T_459 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_496 = _payload_T_462 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_497 = _payload_T_467 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_498 = _payload_T_472 ? _payload_T_17 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_499 = _payload_T_477 ? _payload_T_22 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_500 = _payload_T_482 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_501 = _payload_T_487 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_502 = _payload_T_492 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_503 = _payload_T_495 | _payload_T_496; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_504 = _payload_T_503 | _payload_T_497; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_505 = _payload_T_504 | _payload_T_498; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_506 = _payload_T_505 | _payload_T_499; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_507 = _payload_T_506 | _payload_T_500; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_508 = _payload_T_507 | _payload_T_501; // @[Mux.scala 27:73]
  wire [33:0] payload_9 = _payload_T_508 | _payload_T_502; // @[Mux.scala 27:73]
  wire  tree_18_0_9 = payload_9[0]; // @[Mul.scala 384:26]
  wire  tree_19_0_9 = payload_9[1]; // @[Mul.scala 384:26]
  wire  tree_20_0_9 = payload_9[2]; // @[Mul.scala 384:26]
  wire  tree_21_0_9 = payload_9[3]; // @[Mul.scala 384:26]
  wire  tree_22_0_9 = payload_9[4]; // @[Mul.scala 384:26]
  wire  tree_23_0_9 = payload_9[5]; // @[Mul.scala 384:26]
  wire  tree_24_0_9 = payload_9[6]; // @[Mul.scala 384:26]
  wire  tree_25_0_9 = payload_9[7]; // @[Mul.scala 384:26]
  wire  tree_26_0_9 = payload_9[8]; // @[Mul.scala 384:26]
  wire  tree_27_0_9 = payload_9[9]; // @[Mul.scala 384:26]
  wire  tree_28_0_9 = payload_9[10]; // @[Mul.scala 384:26]
  wire  tree_29_0_9 = payload_9[11]; // @[Mul.scala 384:26]
  wire  tree_30_0_9 = payload_9[12]; // @[Mul.scala 384:26]
  wire  tree_31_0_9 = payload_9[13]; // @[Mul.scala 384:26]
  wire  tree_32_0_9 = payload_9[14]; // @[Mul.scala 384:26]
  wire  tree_33_0_9 = payload_9[15]; // @[Mul.scala 384:26]
  wire  tree_34_0_8 = payload_9[16]; // @[Mul.scala 384:26]
  wire  tree_35_0_8 = payload_9[17]; // @[Mul.scala 384:26]
  wire  tree_36_0_7 = payload_9[18]; // @[Mul.scala 384:26]
  wire  tree_37_0_7 = payload_9[19]; // @[Mul.scala 384:26]
  wire  tree_38_0_6 = payload_9[20]; // @[Mul.scala 384:26]
  wire  tree_39_0_6 = payload_9[21]; // @[Mul.scala 384:26]
  wire  tree_40_0_5 = payload_9[22]; // @[Mul.scala 384:26]
  wire  tree_41_0_5 = payload_9[23]; // @[Mul.scala 384:26]
  wire  tree_42_0_4 = payload_9[24]; // @[Mul.scala 384:26]
  wire  tree_43_0_4 = payload_9[25]; // @[Mul.scala 384:26]
  wire  tree_44_0_3 = payload_9[26]; // @[Mul.scala 384:26]
  wire  tree_45_0_3 = payload_9[27]; // @[Mul.scala 384:26]
  wire  tree_46_0_2 = payload_9[28]; // @[Mul.scala 384:26]
  wire  tree_47_0_2 = payload_9[29]; // @[Mul.scala 384:26]
  wire  tree_48_0_1 = payload_9[30]; // @[Mul.scala 384:26]
  wire  tree_49_0_1 = payload_9[31]; // @[Mul.scala 384:26]
  wire  tree_50_0 = payload_9[32]; // @[Mul.scala 384:26]
  wire  tree_51_0 = payload_9[33]; // @[Mul.scala 384:26]
  wire [2:0] booth4_10 = io_op1[21:19]; // @[Mul.scala 338:131]
  wire  _payload_T_510 = booth4_10 == 3'h0; // @[Mul.scala 341:18]
  wire  _payload_T_513 = booth4_10 == 3'h1; // @[Mul.scala 342:18]
  wire  _payload_T_518 = booth4_10 == 3'h2; // @[Mul.scala 343:18]
  wire  _payload_T_523 = booth4_10 == 3'h3; // @[Mul.scala 344:18]
  wire  _payload_T_528 = booth4_10 == 3'h4; // @[Mul.scala 345:18]
  wire  _payload_T_533 = booth4_10 == 3'h5; // @[Mul.scala 346:18]
  wire  _payload_T_538 = booth4_10 == 3'h6; // @[Mul.scala 347:18]
  wire  _payload_T_543 = booth4_10 == 3'h7; // @[Mul.scala 348:18]
  wire [33:0] _payload_T_546 = _payload_T_510 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_547 = _payload_T_513 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_548 = _payload_T_518 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_549 = _payload_T_523 ? _payload_T_17 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_550 = _payload_T_528 ? _payload_T_22 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_551 = _payload_T_533 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_552 = _payload_T_538 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_553 = _payload_T_543 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_554 = _payload_T_546 | _payload_T_547; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_555 = _payload_T_554 | _payload_T_548; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_556 = _payload_T_555 | _payload_T_549; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_557 = _payload_T_556 | _payload_T_550; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_558 = _payload_T_557 | _payload_T_551; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_559 = _payload_T_558 | _payload_T_552; // @[Mux.scala 27:73]
  wire [33:0] payload_10 = _payload_T_559 | _payload_T_553; // @[Mux.scala 27:73]
  wire  tree_20_0_10 = payload_10[0]; // @[Mul.scala 384:26]
  wire  tree_21_0_10 = payload_10[1]; // @[Mul.scala 384:26]
  wire  tree_22_0_10 = payload_10[2]; // @[Mul.scala 384:26]
  wire  tree_23_0_10 = payload_10[3]; // @[Mul.scala 384:26]
  wire  tree_24_0_10 = payload_10[4]; // @[Mul.scala 384:26]
  wire  tree_25_0_10 = payload_10[5]; // @[Mul.scala 384:26]
  wire  tree_26_0_10 = payload_10[6]; // @[Mul.scala 384:26]
  wire  tree_27_0_10 = payload_10[7]; // @[Mul.scala 384:26]
  wire  tree_28_0_10 = payload_10[8]; // @[Mul.scala 384:26]
  wire  tree_29_0_10 = payload_10[9]; // @[Mul.scala 384:26]
  wire  tree_30_0_10 = payload_10[10]; // @[Mul.scala 384:26]
  wire  tree_31_0_10 = payload_10[11]; // @[Mul.scala 384:26]
  wire  tree_32_0_10 = payload_10[12]; // @[Mul.scala 384:26]
  wire  tree_33_0_10 = payload_10[13]; // @[Mul.scala 384:26]
  wire  tree_34_0_9 = payload_10[14]; // @[Mul.scala 384:26]
  wire  tree_35_0_9 = payload_10[15]; // @[Mul.scala 384:26]
  wire  tree_36_0_8 = payload_10[16]; // @[Mul.scala 384:26]
  wire  tree_37_0_8 = payload_10[17]; // @[Mul.scala 384:26]
  wire  tree_38_0_7 = payload_10[18]; // @[Mul.scala 384:26]
  wire  tree_39_0_7 = payload_10[19]; // @[Mul.scala 384:26]
  wire  tree_40_0_6 = payload_10[20]; // @[Mul.scala 384:26]
  wire  tree_41_0_6 = payload_10[21]; // @[Mul.scala 384:26]
  wire  tree_42_0_5 = payload_10[22]; // @[Mul.scala 384:26]
  wire  tree_43_0_5 = payload_10[23]; // @[Mul.scala 384:26]
  wire  tree_44_0_4 = payload_10[24]; // @[Mul.scala 384:26]
  wire  tree_45_0_4 = payload_10[25]; // @[Mul.scala 384:26]
  wire  tree_46_0_3 = payload_10[26]; // @[Mul.scala 384:26]
  wire  tree_47_0_3 = payload_10[27]; // @[Mul.scala 384:26]
  wire  tree_48_0_2 = payload_10[28]; // @[Mul.scala 384:26]
  wire  tree_49_0_2 = payload_10[29]; // @[Mul.scala 384:26]
  wire  tree_50_0_1 = payload_10[30]; // @[Mul.scala 384:26]
  wire  tree_51_0_1 = payload_10[31]; // @[Mul.scala 384:26]
  wire  tree_52_0 = payload_10[32]; // @[Mul.scala 384:26]
  wire  tree_53_0 = payload_10[33]; // @[Mul.scala 384:26]
  wire [2:0] booth4_11 = io_op1[23:21]; // @[Mul.scala 338:131]
  wire  _payload_T_561 = booth4_11 == 3'h0; // @[Mul.scala 341:18]
  wire  _payload_T_564 = booth4_11 == 3'h1; // @[Mul.scala 342:18]
  wire  _payload_T_569 = booth4_11 == 3'h2; // @[Mul.scala 343:18]
  wire  _payload_T_574 = booth4_11 == 3'h3; // @[Mul.scala 344:18]
  wire  _payload_T_579 = booth4_11 == 3'h4; // @[Mul.scala 345:18]
  wire  _payload_T_584 = booth4_11 == 3'h5; // @[Mul.scala 346:18]
  wire  _payload_T_589 = booth4_11 == 3'h6; // @[Mul.scala 347:18]
  wire  _payload_T_594 = booth4_11 == 3'h7; // @[Mul.scala 348:18]
  wire [33:0] _payload_T_597 = _payload_T_561 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_598 = _payload_T_564 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_599 = _payload_T_569 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_600 = _payload_T_574 ? _payload_T_17 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_601 = _payload_T_579 ? _payload_T_22 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_602 = _payload_T_584 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_603 = _payload_T_589 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_604 = _payload_T_594 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_605 = _payload_T_597 | _payload_T_598; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_606 = _payload_T_605 | _payload_T_599; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_607 = _payload_T_606 | _payload_T_600; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_608 = _payload_T_607 | _payload_T_601; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_609 = _payload_T_608 | _payload_T_602; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_610 = _payload_T_609 | _payload_T_603; // @[Mux.scala 27:73]
  wire [33:0] payload_11 = _payload_T_610 | _payload_T_604; // @[Mux.scala 27:73]
  wire  tree_22_0_11 = payload_11[0]; // @[Mul.scala 384:26]
  wire  tree_23_0_11 = payload_11[1]; // @[Mul.scala 384:26]
  wire  tree_24_0_11 = payload_11[2]; // @[Mul.scala 384:26]
  wire  tree_25_0_11 = payload_11[3]; // @[Mul.scala 384:26]
  wire  tree_26_0_11 = payload_11[4]; // @[Mul.scala 384:26]
  wire  tree_27_0_11 = payload_11[5]; // @[Mul.scala 384:26]
  wire  tree_28_0_11 = payload_11[6]; // @[Mul.scala 384:26]
  wire  tree_29_0_11 = payload_11[7]; // @[Mul.scala 384:26]
  wire  tree_30_0_11 = payload_11[8]; // @[Mul.scala 384:26]
  wire  tree_31_0_11 = payload_11[9]; // @[Mul.scala 384:26]
  wire  tree_32_0_11 = payload_11[10]; // @[Mul.scala 384:26]
  wire  tree_33_0_11 = payload_11[11]; // @[Mul.scala 384:26]
  wire  tree_34_0_10 = payload_11[12]; // @[Mul.scala 384:26]
  wire  tree_35_0_10 = payload_11[13]; // @[Mul.scala 384:26]
  wire  tree_36_0_9 = payload_11[14]; // @[Mul.scala 384:26]
  wire  tree_37_0_9 = payload_11[15]; // @[Mul.scala 384:26]
  wire  tree_38_0_8 = payload_11[16]; // @[Mul.scala 384:26]
  wire  tree_39_0_8 = payload_11[17]; // @[Mul.scala 384:26]
  wire  tree_40_0_7 = payload_11[18]; // @[Mul.scala 384:26]
  wire  tree_41_0_7 = payload_11[19]; // @[Mul.scala 384:26]
  wire  tree_42_0_6 = payload_11[20]; // @[Mul.scala 384:26]
  wire  tree_43_0_6 = payload_11[21]; // @[Mul.scala 384:26]
  wire  tree_44_0_5 = payload_11[22]; // @[Mul.scala 384:26]
  wire  tree_45_0_5 = payload_11[23]; // @[Mul.scala 384:26]
  wire  tree_46_0_4 = payload_11[24]; // @[Mul.scala 384:26]
  wire  tree_47_0_4 = payload_11[25]; // @[Mul.scala 384:26]
  wire  tree_48_0_3 = payload_11[26]; // @[Mul.scala 384:26]
  wire  tree_49_0_3 = payload_11[27]; // @[Mul.scala 384:26]
  wire  tree_50_0_2 = payload_11[28]; // @[Mul.scala 384:26]
  wire  tree_51_0_2 = payload_11[29]; // @[Mul.scala 384:26]
  wire  tree_52_0_1 = payload_11[30]; // @[Mul.scala 384:26]
  wire  tree_53_0_1 = payload_11[31]; // @[Mul.scala 384:26]
  wire  tree_54_0 = payload_11[32]; // @[Mul.scala 384:26]
  wire  tree_55_0 = payload_11[33]; // @[Mul.scala 384:26]
  wire [2:0] booth4_12 = io_op1[25:23]; // @[Mul.scala 338:131]
  wire  _payload_T_612 = booth4_12 == 3'h0; // @[Mul.scala 341:18]
  wire  _payload_T_615 = booth4_12 == 3'h1; // @[Mul.scala 342:18]
  wire  _payload_T_620 = booth4_12 == 3'h2; // @[Mul.scala 343:18]
  wire  _payload_T_625 = booth4_12 == 3'h3; // @[Mul.scala 344:18]
  wire  _payload_T_630 = booth4_12 == 3'h4; // @[Mul.scala 345:18]
  wire  _payload_T_635 = booth4_12 == 3'h5; // @[Mul.scala 346:18]
  wire  _payload_T_640 = booth4_12 == 3'h6; // @[Mul.scala 347:18]
  wire  _payload_T_645 = booth4_12 == 3'h7; // @[Mul.scala 348:18]
  wire [33:0] _payload_T_648 = _payload_T_612 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_649 = _payload_T_615 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_650 = _payload_T_620 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_651 = _payload_T_625 ? _payload_T_17 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_652 = _payload_T_630 ? _payload_T_22 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_653 = _payload_T_635 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_654 = _payload_T_640 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_655 = _payload_T_645 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_656 = _payload_T_648 | _payload_T_649; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_657 = _payload_T_656 | _payload_T_650; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_658 = _payload_T_657 | _payload_T_651; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_659 = _payload_T_658 | _payload_T_652; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_660 = _payload_T_659 | _payload_T_653; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_661 = _payload_T_660 | _payload_T_654; // @[Mux.scala 27:73]
  wire [33:0] payload_12 = _payload_T_661 | _payload_T_655; // @[Mux.scala 27:73]
  wire  tree_24_0_12 = payload_12[0]; // @[Mul.scala 384:26]
  wire  tree_25_0_12 = payload_12[1]; // @[Mul.scala 384:26]
  wire  tree_26_0_12 = payload_12[2]; // @[Mul.scala 384:26]
  wire  tree_27_0_12 = payload_12[3]; // @[Mul.scala 384:26]
  wire  tree_28_0_12 = payload_12[4]; // @[Mul.scala 384:26]
  wire  tree_29_0_12 = payload_12[5]; // @[Mul.scala 384:26]
  wire  tree_30_0_12 = payload_12[6]; // @[Mul.scala 384:26]
  wire  tree_31_0_12 = payload_12[7]; // @[Mul.scala 384:26]
  wire  tree_32_0_12 = payload_12[8]; // @[Mul.scala 384:26]
  wire  tree_33_0_12 = payload_12[9]; // @[Mul.scala 384:26]
  wire  tree_34_0_11 = payload_12[10]; // @[Mul.scala 384:26]
  wire  tree_35_0_11 = payload_12[11]; // @[Mul.scala 384:26]
  wire  tree_36_0_10 = payload_12[12]; // @[Mul.scala 384:26]
  wire  tree_37_0_10 = payload_12[13]; // @[Mul.scala 384:26]
  wire  tree_38_0_9 = payload_12[14]; // @[Mul.scala 384:26]
  wire  tree_39_0_9 = payload_12[15]; // @[Mul.scala 384:26]
  wire  tree_40_0_8 = payload_12[16]; // @[Mul.scala 384:26]
  wire  tree_41_0_8 = payload_12[17]; // @[Mul.scala 384:26]
  wire  tree_42_0_7 = payload_12[18]; // @[Mul.scala 384:26]
  wire  tree_43_0_7 = payload_12[19]; // @[Mul.scala 384:26]
  wire  tree_44_0_6 = payload_12[20]; // @[Mul.scala 384:26]
  wire  tree_45_0_6 = payload_12[21]; // @[Mul.scala 384:26]
  wire  tree_46_0_5 = payload_12[22]; // @[Mul.scala 384:26]
  wire  tree_47_0_5 = payload_12[23]; // @[Mul.scala 384:26]
  wire  tree_48_0_4 = payload_12[24]; // @[Mul.scala 384:26]
  wire  tree_49_0_4 = payload_12[25]; // @[Mul.scala 384:26]
  wire  tree_50_0_3 = payload_12[26]; // @[Mul.scala 384:26]
  wire  tree_51_0_3 = payload_12[27]; // @[Mul.scala 384:26]
  wire  tree_52_0_2 = payload_12[28]; // @[Mul.scala 384:26]
  wire  tree_53_0_2 = payload_12[29]; // @[Mul.scala 384:26]
  wire  tree_54_0_1 = payload_12[30]; // @[Mul.scala 384:26]
  wire  tree_55_0_1 = payload_12[31]; // @[Mul.scala 384:26]
  wire  tree_56_0 = payload_12[32]; // @[Mul.scala 384:26]
  wire  tree_57_0 = payload_12[33]; // @[Mul.scala 384:26]
  wire [2:0] booth4_13 = io_op1[27:25]; // @[Mul.scala 338:131]
  wire  _payload_T_663 = booth4_13 == 3'h0; // @[Mul.scala 341:18]
  wire  _payload_T_666 = booth4_13 == 3'h1; // @[Mul.scala 342:18]
  wire  _payload_T_671 = booth4_13 == 3'h2; // @[Mul.scala 343:18]
  wire  _payload_T_676 = booth4_13 == 3'h3; // @[Mul.scala 344:18]
  wire  _payload_T_681 = booth4_13 == 3'h4; // @[Mul.scala 345:18]
  wire  _payload_T_686 = booth4_13 == 3'h5; // @[Mul.scala 346:18]
  wire  _payload_T_691 = booth4_13 == 3'h6; // @[Mul.scala 347:18]
  wire  _payload_T_696 = booth4_13 == 3'h7; // @[Mul.scala 348:18]
  wire [33:0] _payload_T_699 = _payload_T_663 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_700 = _payload_T_666 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_701 = _payload_T_671 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_702 = _payload_T_676 ? _payload_T_17 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_703 = _payload_T_681 ? _payload_T_22 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_704 = _payload_T_686 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_705 = _payload_T_691 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_706 = _payload_T_696 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_707 = _payload_T_699 | _payload_T_700; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_708 = _payload_T_707 | _payload_T_701; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_709 = _payload_T_708 | _payload_T_702; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_710 = _payload_T_709 | _payload_T_703; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_711 = _payload_T_710 | _payload_T_704; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_712 = _payload_T_711 | _payload_T_705; // @[Mux.scala 27:73]
  wire [33:0] payload_13 = _payload_T_712 | _payload_T_706; // @[Mux.scala 27:73]
  wire  tree_26_0_13 = payload_13[0]; // @[Mul.scala 384:26]
  wire  tree_27_0_13 = payload_13[1]; // @[Mul.scala 384:26]
  wire  tree_28_0_13 = payload_13[2]; // @[Mul.scala 384:26]
  wire  tree_29_0_13 = payload_13[3]; // @[Mul.scala 384:26]
  wire  tree_30_0_13 = payload_13[4]; // @[Mul.scala 384:26]
  wire  tree_31_0_13 = payload_13[5]; // @[Mul.scala 384:26]
  wire  tree_32_0_13 = payload_13[6]; // @[Mul.scala 384:26]
  wire  tree_33_0_13 = payload_13[7]; // @[Mul.scala 384:26]
  wire  tree_34_0_12 = payload_13[8]; // @[Mul.scala 384:26]
  wire  tree_35_0_12 = payload_13[9]; // @[Mul.scala 384:26]
  wire  tree_36_0_11 = payload_13[10]; // @[Mul.scala 384:26]
  wire  tree_37_0_11 = payload_13[11]; // @[Mul.scala 384:26]
  wire  tree_38_0_10 = payload_13[12]; // @[Mul.scala 384:26]
  wire  tree_39_0_10 = payload_13[13]; // @[Mul.scala 384:26]
  wire  tree_40_0_9 = payload_13[14]; // @[Mul.scala 384:26]
  wire  tree_41_0_9 = payload_13[15]; // @[Mul.scala 384:26]
  wire  tree_42_0_8 = payload_13[16]; // @[Mul.scala 384:26]
  wire  tree_43_0_8 = payload_13[17]; // @[Mul.scala 384:26]
  wire  tree_44_0_7 = payload_13[18]; // @[Mul.scala 384:26]
  wire  tree_45_0_7 = payload_13[19]; // @[Mul.scala 384:26]
  wire  tree_46_0_6 = payload_13[20]; // @[Mul.scala 384:26]
  wire  tree_47_0_6 = payload_13[21]; // @[Mul.scala 384:26]
  wire  tree_48_0_5 = payload_13[22]; // @[Mul.scala 384:26]
  wire  tree_49_0_5 = payload_13[23]; // @[Mul.scala 384:26]
  wire  tree_50_0_4 = payload_13[24]; // @[Mul.scala 384:26]
  wire  tree_51_0_4 = payload_13[25]; // @[Mul.scala 384:26]
  wire  tree_52_0_3 = payload_13[26]; // @[Mul.scala 384:26]
  wire  tree_53_0_3 = payload_13[27]; // @[Mul.scala 384:26]
  wire  tree_54_0_2 = payload_13[28]; // @[Mul.scala 384:26]
  wire  tree_55_0_2 = payload_13[29]; // @[Mul.scala 384:26]
  wire  tree_56_0_1 = payload_13[30]; // @[Mul.scala 384:26]
  wire  tree_57_0_1 = payload_13[31]; // @[Mul.scala 384:26]
  wire  tree_58_0 = payload_13[32]; // @[Mul.scala 384:26]
  wire  tree_59_0 = payload_13[33]; // @[Mul.scala 384:26]
  wire [2:0] booth4_14 = io_op1[29:27]; // @[Mul.scala 338:131]
  wire  _payload_T_714 = booth4_14 == 3'h0; // @[Mul.scala 341:18]
  wire  _payload_T_717 = booth4_14 == 3'h1; // @[Mul.scala 342:18]
  wire  _payload_T_722 = booth4_14 == 3'h2; // @[Mul.scala 343:18]
  wire  _payload_T_727 = booth4_14 == 3'h3; // @[Mul.scala 344:18]
  wire  _payload_T_732 = booth4_14 == 3'h4; // @[Mul.scala 345:18]
  wire  _payload_T_737 = booth4_14 == 3'h5; // @[Mul.scala 346:18]
  wire  _payload_T_742 = booth4_14 == 3'h6; // @[Mul.scala 347:18]
  wire  _payload_T_747 = booth4_14 == 3'h7; // @[Mul.scala 348:18]
  wire [33:0] _payload_T_750 = _payload_T_714 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_751 = _payload_T_717 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_752 = _payload_T_722 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_753 = _payload_T_727 ? _payload_T_17 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_754 = _payload_T_732 ? _payload_T_22 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_755 = _payload_T_737 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_756 = _payload_T_742 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_757 = _payload_T_747 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_758 = _payload_T_750 | _payload_T_751; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_759 = _payload_T_758 | _payload_T_752; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_760 = _payload_T_759 | _payload_T_753; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_761 = _payload_T_760 | _payload_T_754; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_762 = _payload_T_761 | _payload_T_755; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_763 = _payload_T_762 | _payload_T_756; // @[Mux.scala 27:73]
  wire [33:0] payload_14 = _payload_T_763 | _payload_T_757; // @[Mux.scala 27:73]
  wire  tree_28_0_14 = payload_14[0]; // @[Mul.scala 384:26]
  wire  tree_29_0_14 = payload_14[1]; // @[Mul.scala 384:26]
  wire  tree_30_0_14 = payload_14[2]; // @[Mul.scala 384:26]
  wire  tree_31_0_14 = payload_14[3]; // @[Mul.scala 384:26]
  wire  tree_32_0_14 = payload_14[4]; // @[Mul.scala 384:26]
  wire  tree_33_0_14 = payload_14[5]; // @[Mul.scala 384:26]
  wire  tree_34_0_13 = payload_14[6]; // @[Mul.scala 384:26]
  wire  tree_35_0_13 = payload_14[7]; // @[Mul.scala 384:26]
  wire  tree_36_0_12 = payload_14[8]; // @[Mul.scala 384:26]
  wire  tree_37_0_12 = payload_14[9]; // @[Mul.scala 384:26]
  wire  tree_38_0_11 = payload_14[10]; // @[Mul.scala 384:26]
  wire  tree_39_0_11 = payload_14[11]; // @[Mul.scala 384:26]
  wire  tree_40_0_10 = payload_14[12]; // @[Mul.scala 384:26]
  wire  tree_41_0_10 = payload_14[13]; // @[Mul.scala 384:26]
  wire  tree_42_0_9 = payload_14[14]; // @[Mul.scala 384:26]
  wire  tree_43_0_9 = payload_14[15]; // @[Mul.scala 384:26]
  wire  tree_44_0_8 = payload_14[16]; // @[Mul.scala 384:26]
  wire  tree_45_0_8 = payload_14[17]; // @[Mul.scala 384:26]
  wire  tree_46_0_7 = payload_14[18]; // @[Mul.scala 384:26]
  wire  tree_47_0_7 = payload_14[19]; // @[Mul.scala 384:26]
  wire  tree_48_0_6 = payload_14[20]; // @[Mul.scala 384:26]
  wire  tree_49_0_6 = payload_14[21]; // @[Mul.scala 384:26]
  wire  tree_50_0_5 = payload_14[22]; // @[Mul.scala 384:26]
  wire  tree_51_0_5 = payload_14[23]; // @[Mul.scala 384:26]
  wire  tree_52_0_4 = payload_14[24]; // @[Mul.scala 384:26]
  wire  tree_53_0_4 = payload_14[25]; // @[Mul.scala 384:26]
  wire  tree_54_0_3 = payload_14[26]; // @[Mul.scala 384:26]
  wire  tree_55_0_3 = payload_14[27]; // @[Mul.scala 384:26]
  wire  tree_56_0_2 = payload_14[28]; // @[Mul.scala 384:26]
  wire  tree_57_0_2 = payload_14[29]; // @[Mul.scala 384:26]
  wire  tree_58_0_1 = payload_14[30]; // @[Mul.scala 384:26]
  wire  tree_59_0_1 = payload_14[31]; // @[Mul.scala 384:26]
  wire  tree_60_0 = payload_14[32]; // @[Mul.scala 384:26]
  wire  tree_61_0 = payload_14[33]; // @[Mul.scala 384:26]
  wire [2:0] booth4_15 = io_op1[31:29]; // @[Mul.scala 338:131]
  wire  _payload_T_765 = booth4_15 == 3'h0; // @[Mul.scala 341:18]
  wire  _payload_T_768 = booth4_15 == 3'h1; // @[Mul.scala 342:18]
  wire  _payload_T_773 = booth4_15 == 3'h2; // @[Mul.scala 343:18]
  wire  _payload_T_778 = booth4_15 == 3'h3; // @[Mul.scala 344:18]
  wire  _payload_T_783 = booth4_15 == 3'h4; // @[Mul.scala 345:18]
  wire  _payload_T_788 = booth4_15 == 3'h5; // @[Mul.scala 346:18]
  wire  _payload_T_793 = booth4_15 == 3'h6; // @[Mul.scala 347:18]
  wire  _payload_T_798 = booth4_15 == 3'h7; // @[Mul.scala 348:18]
  wire [33:0] _payload_T_801 = _payload_T_765 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_802 = _payload_T_768 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_803 = _payload_T_773 ? _payload_T_7 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_804 = _payload_T_778 ? _payload_T_17 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_805 = _payload_T_783 ? _payload_T_22 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_806 = _payload_T_788 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_807 = _payload_T_793 ? _payload_T_27 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_808 = _payload_T_798 ? 34'h300000000 : 34'h0; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_809 = _payload_T_801 | _payload_T_802; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_810 = _payload_T_809 | _payload_T_803; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_811 = _payload_T_810 | _payload_T_804; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_812 = _payload_T_811 | _payload_T_805; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_813 = _payload_T_812 | _payload_T_806; // @[Mux.scala 27:73]
  wire [33:0] _payload_T_814 = _payload_T_813 | _payload_T_807; // @[Mux.scala 27:73]
  wire [33:0] payload_15 = _payload_T_814 | _payload_T_808; // @[Mux.scala 27:73]
  wire  tree_30_0_15 = payload_15[0]; // @[Mul.scala 384:26]
  wire  tree_31_0_15 = payload_15[1]; // @[Mul.scala 384:26]
  wire  tree_32_0_15 = payload_15[2]; // @[Mul.scala 384:26]
  wire  tree_33_0_15 = payload_15[3]; // @[Mul.scala 384:26]
  wire  tree_34_0_14 = payload_15[4]; // @[Mul.scala 384:26]
  wire  tree_35_0_14 = payload_15[5]; // @[Mul.scala 384:26]
  wire  tree_36_0_13 = payload_15[6]; // @[Mul.scala 384:26]
  wire  tree_37_0_13 = payload_15[7]; // @[Mul.scala 384:26]
  wire  tree_38_0_12 = payload_15[8]; // @[Mul.scala 384:26]
  wire  tree_39_0_12 = payload_15[9]; // @[Mul.scala 384:26]
  wire  tree_40_0_11 = payload_15[10]; // @[Mul.scala 384:26]
  wire  tree_41_0_11 = payload_15[11]; // @[Mul.scala 384:26]
  wire  tree_42_0_10 = payload_15[12]; // @[Mul.scala 384:26]
  wire  tree_43_0_10 = payload_15[13]; // @[Mul.scala 384:26]
  wire  tree_44_0_9 = payload_15[14]; // @[Mul.scala 384:26]
  wire  tree_45_0_9 = payload_15[15]; // @[Mul.scala 384:26]
  wire  tree_46_0_8 = payload_15[16]; // @[Mul.scala 384:26]
  wire  tree_47_0_8 = payload_15[17]; // @[Mul.scala 384:26]
  wire  tree_48_0_7 = payload_15[18]; // @[Mul.scala 384:26]
  wire  tree_49_0_7 = payload_15[19]; // @[Mul.scala 384:26]
  wire  tree_50_0_6 = payload_15[20]; // @[Mul.scala 384:26]
  wire  tree_51_0_6 = payload_15[21]; // @[Mul.scala 384:26]
  wire  tree_52_0_5 = payload_15[22]; // @[Mul.scala 384:26]
  wire  tree_53_0_5 = payload_15[23]; // @[Mul.scala 384:26]
  wire  tree_54_0_4 = payload_15[24]; // @[Mul.scala 384:26]
  wire  tree_55_0_4 = payload_15[25]; // @[Mul.scala 384:26]
  wire  tree_56_0_3 = payload_15[26]; // @[Mul.scala 384:26]
  wire  tree_57_0_3 = payload_15[27]; // @[Mul.scala 384:26]
  wire  tree_58_0_2 = payload_15[28]; // @[Mul.scala 384:26]
  wire  tree_59_0_2 = payload_15[29]; // @[Mul.scala 384:26]
  wire  tree_60_0_1 = payload_15[30]; // @[Mul.scala 384:26]
  wire  tree_61_0_1 = payload_15[31]; // @[Mul.scala 384:26]
  wire  tree_62_0 = payload_15[32]; // @[Mul.scala 384:26]
  wire  tree_63_0 = payload_15[33]; // @[Mul.scala 384:26]
  wire  sum = tree_2_0 ^ tree_2_0_1; // @[Mul.scala 206:34]
  wire  cout = tree_2_0 & tree_2_0_1; // @[Mul.scala 207:34]
  wire  sum_1 = tree_3_0 ^ tree_3_0_1; // @[Mul.scala 206:34]
  wire  cout_1 = tree_3_0 & tree_3_0_1; // @[Mul.scala 207:34]
  wire  _sum_T_2 = tree_4_0 ^ tree_4_0_1; // @[Mul.scala 191:34]
  wire  sum_2 = tree_4_0 ^ tree_4_0_1 ^ tree_4_0_2; // @[Mul.scala 191:42]
  wire  cout_2 = tree_4_0 & tree_4_0_1 | _sum_T_2 & tree_4_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_4 = tree_5_0 ^ tree_5_0_1; // @[Mul.scala 191:34]
  wire  sum_3 = tree_5_0 ^ tree_5_0_1 ^ tree_5_0_2; // @[Mul.scala 191:42]
  wire  cout_3 = tree_5_0 & tree_5_0_1 | _sum_T_4 & tree_5_0_2; // @[Mul.scala 192:44]
  wire  sum_4 = tree_6_0 ^ tree_6_0_1; // @[Mul.scala 206:34]
  wire  cout_4 = tree_6_0 & tree_6_0_1; // @[Mul.scala 207:34]
  wire  sum_5 = tree_6_0_2 ^ tree_6_0_3; // @[Mul.scala 206:34]
  wire  cout_5 = tree_6_0_2 & tree_6_0_3; // @[Mul.scala 207:34]
  wire  sum_6 = tree_7_0 ^ tree_7_0_1; // @[Mul.scala 206:34]
  wire  cout_6 = tree_7_0 & tree_7_0_1; // @[Mul.scala 207:34]
  wire  sum_7 = tree_7_0_2 ^ tree_7_0_3; // @[Mul.scala 206:34]
  wire  cout_7 = tree_7_0_2 & tree_7_0_3; // @[Mul.scala 207:34]
  wire  _sum_T_10 = tree_8_0 ^ tree_8_0_1; // @[Mul.scala 191:34]
  wire  sum_8 = tree_8_0 ^ tree_8_0_1 ^ tree_8_0_2; // @[Mul.scala 191:42]
  wire  cout_8 = tree_8_0 & tree_8_0_1 | _sum_T_10 & tree_8_0_2; // @[Mul.scala 192:44]
  wire  ssum_0 = tree_8_0_3 ^ tree_8_0_4; // @[Mul.scala 206:34]
  wire  scout_0 = tree_8_0_3 & tree_8_0_4; // @[Mul.scala 207:34]
  wire  _sum_T_13 = tree_9_0 ^ tree_9_0_1; // @[Mul.scala 191:34]
  wire  sum_9 = tree_9_0 ^ tree_9_0_1 ^ tree_9_0_2; // @[Mul.scala 191:42]
  wire  cout_9 = tree_9_0 & tree_9_0_1 | _sum_T_13 & tree_9_0_2; // @[Mul.scala 192:44]
  wire  ssum_0_1 = tree_9_0_3 ^ tree_9_0_4; // @[Mul.scala 206:34]
  wire  scout_0_1 = tree_9_0_3 & tree_9_0_4; // @[Mul.scala 207:34]
  wire  _sum_T_16 = tree_10_0 ^ tree_10_0_1; // @[Mul.scala 191:34]
  wire  sum_10 = tree_10_0 ^ tree_10_0_1 ^ tree_10_0_2; // @[Mul.scala 191:42]
  wire  cout_10 = tree_10_0 & tree_10_0_1 | _sum_T_16 & tree_10_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_18 = tree_10_0_3 ^ tree_10_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_2 = tree_10_0_3 ^ tree_10_0_4 ^ tree_10_0_5; // @[Mul.scala 191:42]
  wire  scout_0_2 = tree_10_0_3 & tree_10_0_4 | _sum_T_18 & tree_10_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_20 = tree_11_0 ^ tree_11_0_1; // @[Mul.scala 191:34]
  wire  sum_11 = tree_11_0 ^ tree_11_0_1 ^ tree_11_0_2; // @[Mul.scala 191:42]
  wire  cout_11 = tree_11_0 & tree_11_0_1 | _sum_T_20 & tree_11_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_22 = tree_11_0_3 ^ tree_11_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_3 = tree_11_0_3 ^ tree_11_0_4 ^ tree_11_0_5; // @[Mul.scala 191:42]
  wire  scout_0_3 = tree_11_0_3 & tree_11_0_4 | _sum_T_22 & tree_11_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_24 = tree_12_0 ^ tree_12_0_1; // @[Mul.scala 191:34]
  wire  sum_12 = tree_12_0 ^ tree_12_0_1 ^ tree_12_0_2; // @[Mul.scala 191:42]
  wire  cout_12 = tree_12_0 & tree_12_0_1 | _sum_T_24 & tree_12_0_2; // @[Mul.scala 192:44]
  wire  ssum_0_4 = tree_12_0_3 ^ tree_12_0_4; // @[Mul.scala 206:34]
  wire  scout_0_4 = tree_12_0_3 & tree_12_0_4; // @[Mul.scala 207:34]
  wire  ssum_1 = tree_12_0_5 ^ tree_12_0_6; // @[Mul.scala 206:34]
  wire  scout_1 = tree_12_0_5 & tree_12_0_6; // @[Mul.scala 207:34]
  wire  _sum_T_28 = tree_13_0 ^ tree_13_0_1; // @[Mul.scala 191:34]
  wire  sum_13 = tree_13_0 ^ tree_13_0_1 ^ tree_13_0_2; // @[Mul.scala 191:42]
  wire  cout_13 = tree_13_0 & tree_13_0_1 | _sum_T_28 & tree_13_0_2; // @[Mul.scala 192:44]
  wire  ssum_0_5 = tree_13_0_3 ^ tree_13_0_4; // @[Mul.scala 206:34]
  wire  scout_0_5 = tree_13_0_3 & tree_13_0_4; // @[Mul.scala 207:34]
  wire  ssum_1_1 = tree_13_0_5 ^ tree_13_0_6; // @[Mul.scala 206:34]
  wire  scout_1_1 = tree_13_0_5 & tree_13_0_6; // @[Mul.scala 207:34]
  wire  _sum_T_32 = tree_14_0 ^ tree_14_0_1; // @[Mul.scala 191:34]
  wire  sum_14 = tree_14_0 ^ tree_14_0_1 ^ tree_14_0_2; // @[Mul.scala 191:42]
  wire  cout_14 = tree_14_0 & tree_14_0_1 | _sum_T_32 & tree_14_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_34 = tree_14_0_3 ^ tree_14_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_6 = tree_14_0_3 ^ tree_14_0_4 ^ tree_14_0_5; // @[Mul.scala 191:42]
  wire  scout_0_6 = tree_14_0_3 & tree_14_0_4 | _sum_T_34 & tree_14_0_5; // @[Mul.scala 192:44]
  wire  ssum_1_2 = tree_14_0_6 ^ tree_14_0_7; // @[Mul.scala 206:34]
  wire  scout_1_2 = tree_14_0_6 & tree_14_0_7; // @[Mul.scala 207:34]
  wire  _sum_T_37 = tree_15_0 ^ tree_15_0_1; // @[Mul.scala 191:34]
  wire  sum_15 = tree_15_0 ^ tree_15_0_1 ^ tree_15_0_2; // @[Mul.scala 191:42]
  wire  cout_15 = tree_15_0 & tree_15_0_1 | _sum_T_37 & tree_15_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_39 = tree_15_0_3 ^ tree_15_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_7 = tree_15_0_3 ^ tree_15_0_4 ^ tree_15_0_5; // @[Mul.scala 191:42]
  wire  scout_0_7 = tree_15_0_3 & tree_15_0_4 | _sum_T_39 & tree_15_0_5; // @[Mul.scala 192:44]
  wire  ssum_1_3 = tree_15_0_6 ^ tree_15_0_7; // @[Mul.scala 206:34]
  wire  scout_1_3 = tree_15_0_6 & tree_15_0_7; // @[Mul.scala 207:34]
  wire  _sum_T_42 = tree_16_0 ^ tree_16_0_1; // @[Mul.scala 191:34]
  wire  sum_16 = tree_16_0 ^ tree_16_0_1 ^ tree_16_0_2; // @[Mul.scala 191:42]
  wire  cout_16 = tree_16_0 & tree_16_0_1 | _sum_T_42 & tree_16_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_44 = tree_16_0_3 ^ tree_16_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_8 = tree_16_0_3 ^ tree_16_0_4 ^ tree_16_0_5; // @[Mul.scala 191:42]
  wire  scout_0_8 = tree_16_0_3 & tree_16_0_4 | _sum_T_44 & tree_16_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_46 = tree_16_0_6 ^ tree_16_0_7; // @[Mul.scala 191:34]
  wire  ssum_1_4 = tree_16_0_6 ^ tree_16_0_7 ^ tree_16_0_8; // @[Mul.scala 191:42]
  wire  scout_1_4 = tree_16_0_6 & tree_16_0_7 | _sum_T_46 & tree_16_0_8; // @[Mul.scala 192:44]
  wire  _sum_T_48 = tree_17_0 ^ tree_17_0_1; // @[Mul.scala 191:34]
  wire  sum_17 = tree_17_0 ^ tree_17_0_1 ^ tree_17_0_2; // @[Mul.scala 191:42]
  wire  cout_17 = tree_17_0 & tree_17_0_1 | _sum_T_48 & tree_17_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_50 = tree_17_0_3 ^ tree_17_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_9 = tree_17_0_3 ^ tree_17_0_4 ^ tree_17_0_5; // @[Mul.scala 191:42]
  wire  scout_0_9 = tree_17_0_3 & tree_17_0_4 | _sum_T_50 & tree_17_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_52 = tree_17_0_6 ^ tree_17_0_7; // @[Mul.scala 191:34]
  wire  ssum_1_5 = tree_17_0_6 ^ tree_17_0_7 ^ tree_17_0_8; // @[Mul.scala 191:42]
  wire  scout_1_5 = tree_17_0_6 & tree_17_0_7 | _sum_T_52 & tree_17_0_8; // @[Mul.scala 192:44]
  wire  _sum_T_54 = tree_18_0 ^ tree_18_0_1; // @[Mul.scala 191:34]
  wire  sum_18 = tree_18_0 ^ tree_18_0_1 ^ tree_18_0_2; // @[Mul.scala 191:42]
  wire  cout_18 = tree_18_0 & tree_18_0_1 | _sum_T_54 & tree_18_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_56 = tree_18_0_3 ^ tree_18_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_10 = tree_18_0_3 ^ tree_18_0_4 ^ tree_18_0_5; // @[Mul.scala 191:42]
  wire  scout_0_10 = tree_18_0_3 & tree_18_0_4 | _sum_T_56 & tree_18_0_5; // @[Mul.scala 192:44]
  wire  ssum_1_6 = tree_18_0_6 ^ tree_18_0_7; // @[Mul.scala 206:34]
  wire  scout_1_6 = tree_18_0_6 & tree_18_0_7; // @[Mul.scala 207:34]
  wire  ssum_2 = tree_18_0_8 ^ tree_18_0_9; // @[Mul.scala 206:34]
  wire  scout_2 = tree_18_0_8 & tree_18_0_9; // @[Mul.scala 207:34]
  wire  _sum_T_60 = tree_19_0 ^ tree_19_0_1; // @[Mul.scala 191:34]
  wire  sum_19 = tree_19_0 ^ tree_19_0_1 ^ tree_19_0_2; // @[Mul.scala 191:42]
  wire  cout_19 = tree_19_0 & tree_19_0_1 | _sum_T_60 & tree_19_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_62 = tree_19_0_3 ^ tree_19_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_11 = tree_19_0_3 ^ tree_19_0_4 ^ tree_19_0_5; // @[Mul.scala 191:42]
  wire  scout_0_11 = tree_19_0_3 & tree_19_0_4 | _sum_T_62 & tree_19_0_5; // @[Mul.scala 192:44]
  wire  ssum_1_7 = tree_19_0_6 ^ tree_19_0_7; // @[Mul.scala 206:34]
  wire  scout_1_7 = tree_19_0_6 & tree_19_0_7; // @[Mul.scala 207:34]
  wire  ssum_2_1 = tree_19_0_8 ^ tree_19_0_9; // @[Mul.scala 206:34]
  wire  scout_2_1 = tree_19_0_8 & tree_19_0_9; // @[Mul.scala 207:34]
  wire  _sum_T_66 = tree_20_0 ^ tree_20_0_1; // @[Mul.scala 191:34]
  wire  sum_20 = tree_20_0 ^ tree_20_0_1 ^ tree_20_0_2; // @[Mul.scala 191:42]
  wire  cout_20 = tree_20_0 & tree_20_0_1 | _sum_T_66 & tree_20_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_68 = tree_20_0_3 ^ tree_20_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_12 = tree_20_0_3 ^ tree_20_0_4 ^ tree_20_0_5; // @[Mul.scala 191:42]
  wire  scout_0_12 = tree_20_0_3 & tree_20_0_4 | _sum_T_68 & tree_20_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_70 = tree_20_0_6 ^ tree_20_0_7; // @[Mul.scala 191:34]
  wire  ssum_1_8 = tree_20_0_6 ^ tree_20_0_7 ^ tree_20_0_8; // @[Mul.scala 191:42]
  wire  scout_1_8 = tree_20_0_6 & tree_20_0_7 | _sum_T_70 & tree_20_0_8; // @[Mul.scala 192:44]
  wire  ssum_2_2 = tree_20_0_9 ^ tree_20_0_10; // @[Mul.scala 206:34]
  wire  scout_2_2 = tree_20_0_9 & tree_20_0_10; // @[Mul.scala 207:34]
  wire  _sum_T_73 = tree_21_0 ^ tree_21_0_1; // @[Mul.scala 191:34]
  wire  sum_21 = tree_21_0 ^ tree_21_0_1 ^ tree_21_0_2; // @[Mul.scala 191:42]
  wire  cout_21 = tree_21_0 & tree_21_0_1 | _sum_T_73 & tree_21_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_75 = tree_21_0_3 ^ tree_21_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_13 = tree_21_0_3 ^ tree_21_0_4 ^ tree_21_0_5; // @[Mul.scala 191:42]
  wire  scout_0_13 = tree_21_0_3 & tree_21_0_4 | _sum_T_75 & tree_21_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_77 = tree_21_0_6 ^ tree_21_0_7; // @[Mul.scala 191:34]
  wire  ssum_1_9 = tree_21_0_6 ^ tree_21_0_7 ^ tree_21_0_8; // @[Mul.scala 191:42]
  wire  scout_1_9 = tree_21_0_6 & tree_21_0_7 | _sum_T_77 & tree_21_0_8; // @[Mul.scala 192:44]
  wire  ssum_2_3 = tree_21_0_9 ^ tree_21_0_10; // @[Mul.scala 206:34]
  wire  scout_2_3 = tree_21_0_9 & tree_21_0_10; // @[Mul.scala 207:34]
  wire  _sum_T_80 = tree_22_0 ^ tree_22_0_1; // @[Mul.scala 191:34]
  wire  sum_22 = tree_22_0 ^ tree_22_0_1 ^ tree_22_0_2; // @[Mul.scala 191:42]
  wire  cout_22 = tree_22_0 & tree_22_0_1 | _sum_T_80 & tree_22_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_82 = tree_22_0_3 ^ tree_22_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_14 = tree_22_0_3 ^ tree_22_0_4 ^ tree_22_0_5; // @[Mul.scala 191:42]
  wire  scout_0_14 = tree_22_0_3 & tree_22_0_4 | _sum_T_82 & tree_22_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_84 = tree_22_0_6 ^ tree_22_0_7; // @[Mul.scala 191:34]
  wire  ssum_1_10 = tree_22_0_6 ^ tree_22_0_7 ^ tree_22_0_8; // @[Mul.scala 191:42]
  wire  scout_1_10 = tree_22_0_6 & tree_22_0_7 | _sum_T_84 & tree_22_0_8; // @[Mul.scala 192:44]
  wire  _sum_T_86 = tree_22_0_9 ^ tree_22_0_10; // @[Mul.scala 191:34]
  wire  ssum_2_4 = tree_22_0_9 ^ tree_22_0_10 ^ tree_22_0_11; // @[Mul.scala 191:42]
  wire  scout_2_4 = tree_22_0_9 & tree_22_0_10 | _sum_T_86 & tree_22_0_11; // @[Mul.scala 192:44]
  wire  _sum_T_88 = tree_23_0 ^ tree_23_0_1; // @[Mul.scala 191:34]
  wire  sum_23 = tree_23_0 ^ tree_23_0_1 ^ tree_23_0_2; // @[Mul.scala 191:42]
  wire  cout_23 = tree_23_0 & tree_23_0_1 | _sum_T_88 & tree_23_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_90 = tree_23_0_3 ^ tree_23_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_15 = tree_23_0_3 ^ tree_23_0_4 ^ tree_23_0_5; // @[Mul.scala 191:42]
  wire  scout_0_15 = tree_23_0_3 & tree_23_0_4 | _sum_T_90 & tree_23_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_92 = tree_23_0_6 ^ tree_23_0_7; // @[Mul.scala 191:34]
  wire  ssum_1_11 = tree_23_0_6 ^ tree_23_0_7 ^ tree_23_0_8; // @[Mul.scala 191:42]
  wire  scout_1_11 = tree_23_0_6 & tree_23_0_7 | _sum_T_92 & tree_23_0_8; // @[Mul.scala 192:44]
  wire  _sum_T_94 = tree_23_0_9 ^ tree_23_0_10; // @[Mul.scala 191:34]
  wire  ssum_2_5 = tree_23_0_9 ^ tree_23_0_10 ^ tree_23_0_11; // @[Mul.scala 191:42]
  wire  scout_2_5 = tree_23_0_9 & tree_23_0_10 | _sum_T_94 & tree_23_0_11; // @[Mul.scala 192:44]
  wire  _sum_T_96 = tree_24_0 ^ tree_24_0_1; // @[Mul.scala 191:34]
  wire  sum_24 = tree_24_0 ^ tree_24_0_1 ^ tree_24_0_2; // @[Mul.scala 191:42]
  wire  cout_24 = tree_24_0 & tree_24_0_1 | _sum_T_96 & tree_24_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_98 = tree_24_0_3 ^ tree_24_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_16 = tree_24_0_3 ^ tree_24_0_4 ^ tree_24_0_5; // @[Mul.scala 191:42]
  wire  scout_0_16 = tree_24_0_3 & tree_24_0_4 | _sum_T_98 & tree_24_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_100 = tree_24_0_6 ^ tree_24_0_7; // @[Mul.scala 191:34]
  wire  ssum_1_12 = tree_24_0_6 ^ tree_24_0_7 ^ tree_24_0_8; // @[Mul.scala 191:42]
  wire  scout_1_12 = tree_24_0_6 & tree_24_0_7 | _sum_T_100 & tree_24_0_8; // @[Mul.scala 192:44]
  wire  ssum_2_6 = tree_24_0_9 ^ tree_24_0_10; // @[Mul.scala 206:34]
  wire  scout_2_6 = tree_24_0_9 & tree_24_0_10; // @[Mul.scala 207:34]
  wire  ssum_3 = tree_24_0_11 ^ tree_24_0_12; // @[Mul.scala 206:34]
  wire  scout_3 = tree_24_0_11 & tree_24_0_12; // @[Mul.scala 207:34]
  wire  _sum_T_104 = tree_25_0 ^ tree_25_0_1; // @[Mul.scala 191:34]
  wire  sum_25 = tree_25_0 ^ tree_25_0_1 ^ tree_25_0_2; // @[Mul.scala 191:42]
  wire  cout_25 = tree_25_0 & tree_25_0_1 | _sum_T_104 & tree_25_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_106 = tree_25_0_3 ^ tree_25_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_17 = tree_25_0_3 ^ tree_25_0_4 ^ tree_25_0_5; // @[Mul.scala 191:42]
  wire  scout_0_17 = tree_25_0_3 & tree_25_0_4 | _sum_T_106 & tree_25_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_108 = tree_25_0_6 ^ tree_25_0_7; // @[Mul.scala 191:34]
  wire  ssum_1_13 = tree_25_0_6 ^ tree_25_0_7 ^ tree_25_0_8; // @[Mul.scala 191:42]
  wire  scout_1_13 = tree_25_0_6 & tree_25_0_7 | _sum_T_108 & tree_25_0_8; // @[Mul.scala 192:44]
  wire  ssum_2_7 = tree_25_0_9 ^ tree_25_0_10; // @[Mul.scala 206:34]
  wire  scout_2_7 = tree_25_0_9 & tree_25_0_10; // @[Mul.scala 207:34]
  wire  ssum_3_1 = tree_25_0_11 ^ tree_25_0_12; // @[Mul.scala 206:34]
  wire  scout_3_1 = tree_25_0_11 & tree_25_0_12; // @[Mul.scala 207:34]
  wire  _sum_T_112 = tree_26_0 ^ tree_26_0_1; // @[Mul.scala 191:34]
  wire  sum_26 = tree_26_0 ^ tree_26_0_1 ^ tree_26_0_2; // @[Mul.scala 191:42]
  wire  cout_26 = tree_26_0 & tree_26_0_1 | _sum_T_112 & tree_26_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_114 = tree_26_0_3 ^ tree_26_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_18 = tree_26_0_3 ^ tree_26_0_4 ^ tree_26_0_5; // @[Mul.scala 191:42]
  wire  scout_0_18 = tree_26_0_3 & tree_26_0_4 | _sum_T_114 & tree_26_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_116 = tree_26_0_6 ^ tree_26_0_7; // @[Mul.scala 191:34]
  wire  ssum_1_14 = tree_26_0_6 ^ tree_26_0_7 ^ tree_26_0_8; // @[Mul.scala 191:42]
  wire  scout_1_14 = tree_26_0_6 & tree_26_0_7 | _sum_T_116 & tree_26_0_8; // @[Mul.scala 192:44]
  wire  _sum_T_118 = tree_26_0_9 ^ tree_26_0_10; // @[Mul.scala 191:34]
  wire  ssum_2_8 = tree_26_0_9 ^ tree_26_0_10 ^ tree_26_0_11; // @[Mul.scala 191:42]
  wire  scout_2_8 = tree_26_0_9 & tree_26_0_10 | _sum_T_118 & tree_26_0_11; // @[Mul.scala 192:44]
  wire  ssum_3_2 = tree_26_0_12 ^ tree_26_0_13; // @[Mul.scala 206:34]
  wire  scout_3_2 = tree_26_0_12 & tree_26_0_13; // @[Mul.scala 207:34]
  wire  _sum_T_121 = tree_27_0 ^ tree_27_0_1; // @[Mul.scala 191:34]
  wire  sum_27 = tree_27_0 ^ tree_27_0_1 ^ tree_27_0_2; // @[Mul.scala 191:42]
  wire  cout_27 = tree_27_0 & tree_27_0_1 | _sum_T_121 & tree_27_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_123 = tree_27_0_3 ^ tree_27_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_19 = tree_27_0_3 ^ tree_27_0_4 ^ tree_27_0_5; // @[Mul.scala 191:42]
  wire  scout_0_19 = tree_27_0_3 & tree_27_0_4 | _sum_T_123 & tree_27_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_125 = tree_27_0_6 ^ tree_27_0_7; // @[Mul.scala 191:34]
  wire  ssum_1_15 = tree_27_0_6 ^ tree_27_0_7 ^ tree_27_0_8; // @[Mul.scala 191:42]
  wire  scout_1_15 = tree_27_0_6 & tree_27_0_7 | _sum_T_125 & tree_27_0_8; // @[Mul.scala 192:44]
  wire  _sum_T_127 = tree_27_0_9 ^ tree_27_0_10; // @[Mul.scala 191:34]
  wire  ssum_2_9 = tree_27_0_9 ^ tree_27_0_10 ^ tree_27_0_11; // @[Mul.scala 191:42]
  wire  scout_2_9 = tree_27_0_9 & tree_27_0_10 | _sum_T_127 & tree_27_0_11; // @[Mul.scala 192:44]
  wire  ssum_3_3 = tree_27_0_12 ^ tree_27_0_13; // @[Mul.scala 206:34]
  wire  scout_3_3 = tree_27_0_12 & tree_27_0_13; // @[Mul.scala 207:34]
  wire  _sum_T_130 = tree_28_0 ^ tree_28_0_1; // @[Mul.scala 191:34]
  wire  sum_28 = tree_28_0 ^ tree_28_0_1 ^ tree_28_0_2; // @[Mul.scala 191:42]
  wire  cout_28 = tree_28_0 & tree_28_0_1 | _sum_T_130 & tree_28_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_132 = tree_28_0_3 ^ tree_28_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_20 = tree_28_0_3 ^ tree_28_0_4 ^ tree_28_0_5; // @[Mul.scala 191:42]
  wire  scout_0_20 = tree_28_0_3 & tree_28_0_4 | _sum_T_132 & tree_28_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_134 = tree_28_0_6 ^ tree_28_0_7; // @[Mul.scala 191:34]
  wire  ssum_1_16 = tree_28_0_6 ^ tree_28_0_7 ^ tree_28_0_8; // @[Mul.scala 191:42]
  wire  scout_1_16 = tree_28_0_6 & tree_28_0_7 | _sum_T_134 & tree_28_0_8; // @[Mul.scala 192:44]
  wire  _sum_T_136 = tree_28_0_9 ^ tree_28_0_10; // @[Mul.scala 191:34]
  wire  ssum_2_10 = tree_28_0_9 ^ tree_28_0_10 ^ tree_28_0_11; // @[Mul.scala 191:42]
  wire  scout_2_10 = tree_28_0_9 & tree_28_0_10 | _sum_T_136 & tree_28_0_11; // @[Mul.scala 192:44]
  wire  _sum_T_138 = tree_28_0_12 ^ tree_28_0_13; // @[Mul.scala 191:34]
  wire  ssum_3_4 = tree_28_0_12 ^ tree_28_0_13 ^ tree_28_0_14; // @[Mul.scala 191:42]
  wire  scout_3_4 = tree_28_0_12 & tree_28_0_13 | _sum_T_138 & tree_28_0_14; // @[Mul.scala 192:44]
  wire  _sum_T_140 = tree_29_0 ^ tree_29_0_1; // @[Mul.scala 191:34]
  wire  sum_29 = tree_29_0 ^ tree_29_0_1 ^ tree_29_0_2; // @[Mul.scala 191:42]
  wire  cout_29 = tree_29_0 & tree_29_0_1 | _sum_T_140 & tree_29_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_142 = tree_29_0_3 ^ tree_29_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_21 = tree_29_0_3 ^ tree_29_0_4 ^ tree_29_0_5; // @[Mul.scala 191:42]
  wire  scout_0_21 = tree_29_0_3 & tree_29_0_4 | _sum_T_142 & tree_29_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_144 = tree_29_0_6 ^ tree_29_0_7; // @[Mul.scala 191:34]
  wire  ssum_1_17 = tree_29_0_6 ^ tree_29_0_7 ^ tree_29_0_8; // @[Mul.scala 191:42]
  wire  scout_1_17 = tree_29_0_6 & tree_29_0_7 | _sum_T_144 & tree_29_0_8; // @[Mul.scala 192:44]
  wire  _sum_T_146 = tree_29_0_9 ^ tree_29_0_10; // @[Mul.scala 191:34]
  wire  ssum_2_11 = tree_29_0_9 ^ tree_29_0_10 ^ tree_29_0_11; // @[Mul.scala 191:42]
  wire  scout_2_11 = tree_29_0_9 & tree_29_0_10 | _sum_T_146 & tree_29_0_11; // @[Mul.scala 192:44]
  wire  _sum_T_148 = tree_29_0_12 ^ tree_29_0_13; // @[Mul.scala 191:34]
  wire  ssum_3_5 = tree_29_0_12 ^ tree_29_0_13 ^ tree_29_0_14; // @[Mul.scala 191:42]
  wire  scout_3_5 = tree_29_0_12 & tree_29_0_13 | _sum_T_148 & tree_29_0_14; // @[Mul.scala 192:44]
  wire  _sum_T_150 = tree_30_0 ^ tree_30_0_1; // @[Mul.scala 191:34]
  wire  sum_30 = tree_30_0 ^ tree_30_0_1 ^ tree_30_0_2; // @[Mul.scala 191:42]
  wire  cout_30 = tree_30_0 & tree_30_0_1 | _sum_T_150 & tree_30_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_152 = tree_30_0_3 ^ tree_30_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_22 = tree_30_0_3 ^ tree_30_0_4 ^ tree_30_0_5; // @[Mul.scala 191:42]
  wire  scout_0_22 = tree_30_0_3 & tree_30_0_4 | _sum_T_152 & tree_30_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_154 = tree_30_0_6 ^ tree_30_0_7; // @[Mul.scala 191:34]
  wire  ssum_1_18 = tree_30_0_6 ^ tree_30_0_7 ^ tree_30_0_8; // @[Mul.scala 191:42]
  wire  scout_1_18 = tree_30_0_6 & tree_30_0_7 | _sum_T_154 & tree_30_0_8; // @[Mul.scala 192:44]
  wire  _sum_T_156 = tree_30_0_9 ^ tree_30_0_10; // @[Mul.scala 191:34]
  wire  ssum_2_12 = tree_30_0_9 ^ tree_30_0_10 ^ tree_30_0_11; // @[Mul.scala 191:42]
  wire  scout_2_12 = tree_30_0_9 & tree_30_0_10 | _sum_T_156 & tree_30_0_11; // @[Mul.scala 192:44]
  wire  ssum_3_6 = tree_30_0_12 ^ tree_30_0_13; // @[Mul.scala 206:34]
  wire  scout_3_6 = tree_30_0_12 & tree_30_0_13; // @[Mul.scala 207:34]
  wire  ssum_4 = tree_30_0_14 ^ tree_30_0_15; // @[Mul.scala 206:34]
  wire  scout_4 = tree_30_0_14 & tree_30_0_15; // @[Mul.scala 207:34]
  wire  _sum_T_160 = tree_31_0 ^ tree_31_0_1; // @[Mul.scala 191:34]
  wire  sum_31 = tree_31_0 ^ tree_31_0_1 ^ tree_31_0_2; // @[Mul.scala 191:42]
  wire  cout_31 = tree_31_0 & tree_31_0_1 | _sum_T_160 & tree_31_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_162 = tree_31_0_3 ^ tree_31_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_23 = tree_31_0_3 ^ tree_31_0_4 ^ tree_31_0_5; // @[Mul.scala 191:42]
  wire  scout_0_23 = tree_31_0_3 & tree_31_0_4 | _sum_T_162 & tree_31_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_164 = tree_31_0_6 ^ tree_31_0_7; // @[Mul.scala 191:34]
  wire  ssum_1_19 = tree_31_0_6 ^ tree_31_0_7 ^ tree_31_0_8; // @[Mul.scala 191:42]
  wire  scout_1_19 = tree_31_0_6 & tree_31_0_7 | _sum_T_164 & tree_31_0_8; // @[Mul.scala 192:44]
  wire  _sum_T_166 = tree_31_0_9 ^ tree_31_0_10; // @[Mul.scala 191:34]
  wire  ssum_2_13 = tree_31_0_9 ^ tree_31_0_10 ^ tree_31_0_11; // @[Mul.scala 191:42]
  wire  scout_2_13 = tree_31_0_9 & tree_31_0_10 | _sum_T_166 & tree_31_0_11; // @[Mul.scala 192:44]
  wire  ssum_3_7 = tree_31_0_12 ^ tree_31_0_13; // @[Mul.scala 206:34]
  wire  scout_3_7 = tree_31_0_12 & tree_31_0_13; // @[Mul.scala 207:34]
  wire  ssum_4_1 = tree_31_0_14 ^ tree_31_0_15; // @[Mul.scala 206:34]
  wire  scout_4_1 = tree_31_0_14 & tree_31_0_15; // @[Mul.scala 207:34]
  wire  _sum_T_170 = tree_32_0 ^ tree_32_0_1; // @[Mul.scala 191:34]
  wire  sum_32 = tree_32_0 ^ tree_32_0_1 ^ tree_32_0_2; // @[Mul.scala 191:42]
  wire  cout_32 = tree_32_0 & tree_32_0_1 | _sum_T_170 & tree_32_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_172 = tree_32_0_3 ^ tree_32_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_24 = tree_32_0_3 ^ tree_32_0_4 ^ tree_32_0_5; // @[Mul.scala 191:42]
  wire  scout_0_24 = tree_32_0_3 & tree_32_0_4 | _sum_T_172 & tree_32_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_174 = tree_32_0_6 ^ tree_32_0_7; // @[Mul.scala 191:34]
  wire  ssum_1_20 = tree_32_0_6 ^ tree_32_0_7 ^ tree_32_0_8; // @[Mul.scala 191:42]
  wire  scout_1_20 = tree_32_0_6 & tree_32_0_7 | _sum_T_174 & tree_32_0_8; // @[Mul.scala 192:44]
  wire  _sum_T_176 = tree_32_0_9 ^ tree_32_0_10; // @[Mul.scala 191:34]
  wire  ssum_2_14 = tree_32_0_9 ^ tree_32_0_10 ^ tree_32_0_11; // @[Mul.scala 191:42]
  wire  scout_2_14 = tree_32_0_9 & tree_32_0_10 | _sum_T_176 & tree_32_0_11; // @[Mul.scala 192:44]
  wire  _sum_T_178 = tree_32_0_12 ^ tree_32_0_13; // @[Mul.scala 191:34]
  wire  ssum_3_8 = tree_32_0_12 ^ tree_32_0_13 ^ tree_32_0_14; // @[Mul.scala 191:42]
  wire  scout_3_8 = tree_32_0_12 & tree_32_0_13 | _sum_T_178 & tree_32_0_14; // @[Mul.scala 192:44]
  wire  ssum_4_2 = tree_32_0_15 ^ 1'h1; // @[Mul.scala 206:34]
  wire  _sum_T_181 = tree_33_0 ^ tree_33_0_1; // @[Mul.scala 191:34]
  wire  sum_33 = tree_33_0 ^ tree_33_0_1 ^ tree_33_0_2; // @[Mul.scala 191:42]
  wire  cout_33 = tree_33_0 & tree_33_0_1 | _sum_T_181 & tree_33_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_183 = tree_33_0_3 ^ tree_33_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_25 = tree_33_0_3 ^ tree_33_0_4 ^ tree_33_0_5; // @[Mul.scala 191:42]
  wire  scout_0_25 = tree_33_0_3 & tree_33_0_4 | _sum_T_183 & tree_33_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_185 = tree_33_0_6 ^ tree_33_0_7; // @[Mul.scala 191:34]
  wire  ssum_1_21 = tree_33_0_6 ^ tree_33_0_7 ^ tree_33_0_8; // @[Mul.scala 191:42]
  wire  scout_1_21 = tree_33_0_6 & tree_33_0_7 | _sum_T_185 & tree_33_0_8; // @[Mul.scala 192:44]
  wire  _sum_T_187 = tree_33_0_9 ^ tree_33_0_10; // @[Mul.scala 191:34]
  wire  ssum_2_15 = tree_33_0_9 ^ tree_33_0_10 ^ tree_33_0_11; // @[Mul.scala 191:42]
  wire  scout_2_15 = tree_33_0_9 & tree_33_0_10 | _sum_T_187 & tree_33_0_11; // @[Mul.scala 192:44]
  wire  ssum_3_9 = tree_33_0_12 ^ tree_33_0_13; // @[Mul.scala 206:34]
  wire  scout_3_9 = tree_33_0_12 & tree_33_0_13; // @[Mul.scala 207:34]
  wire  ssum_4_3 = tree_33_0_14 ^ tree_33_0_15; // @[Mul.scala 206:34]
  wire  scout_4_3 = tree_33_0_14 & tree_33_0_15; // @[Mul.scala 207:34]
  wire  _sum_T_191 = tree_34_0 ^ tree_34_0_1; // @[Mul.scala 191:34]
  wire  sum_34 = tree_34_0 ^ tree_34_0_1 ^ tree_34_0_2; // @[Mul.scala 191:42]
  wire  cout_34 = tree_34_0 & tree_34_0_1 | _sum_T_191 & tree_34_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_193 = tree_34_0_3 ^ tree_34_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_26 = tree_34_0_3 ^ tree_34_0_4 ^ tree_34_0_5; // @[Mul.scala 191:42]
  wire  scout_0_26 = tree_34_0_3 & tree_34_0_4 | _sum_T_193 & tree_34_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_195 = tree_34_0_6 ^ tree_34_0_7; // @[Mul.scala 191:34]
  wire  ssum_1_22 = tree_34_0_6 ^ tree_34_0_7 ^ tree_34_0_8; // @[Mul.scala 191:42]
  wire  scout_1_22 = tree_34_0_6 & tree_34_0_7 | _sum_T_195 & tree_34_0_8; // @[Mul.scala 192:44]
  wire  _sum_T_197 = tree_34_0_9 ^ tree_34_0_10; // @[Mul.scala 191:34]
  wire  ssum_2_16 = tree_34_0_9 ^ tree_34_0_10 ^ tree_34_0_11; // @[Mul.scala 191:42]
  wire  scout_2_16 = tree_34_0_9 & tree_34_0_10 | _sum_T_197 & tree_34_0_11; // @[Mul.scala 192:44]
  wire  _sum_T_199 = tree_34_0_12 ^ tree_34_0_13; // @[Mul.scala 191:34]
  wire  ssum_3_10 = tree_34_0_12 ^ tree_34_0_13 ^ tree_34_0_14; // @[Mul.scala 191:42]
  wire  scout_3_10 = tree_34_0_12 & tree_34_0_13 | _sum_T_199 & tree_34_0_14; // @[Mul.scala 192:44]
  wire  _sum_T_201 = tree_35_0 ^ tree_35_0_1; // @[Mul.scala 191:34]
  wire  sum_35 = tree_35_0 ^ tree_35_0_1 ^ tree_35_0_2; // @[Mul.scala 191:42]
  wire  cout_35 = tree_35_0 & tree_35_0_1 | _sum_T_201 & tree_35_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_203 = tree_35_0_3 ^ tree_35_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_27 = tree_35_0_3 ^ tree_35_0_4 ^ tree_35_0_5; // @[Mul.scala 191:42]
  wire  scout_0_27 = tree_35_0_3 & tree_35_0_4 | _sum_T_203 & tree_35_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_205 = tree_35_0_6 ^ tree_35_0_7; // @[Mul.scala 191:34]
  wire  ssum_1_23 = tree_35_0_6 ^ tree_35_0_7 ^ tree_35_0_8; // @[Mul.scala 191:42]
  wire  scout_1_23 = tree_35_0_6 & tree_35_0_7 | _sum_T_205 & tree_35_0_8; // @[Mul.scala 192:44]
  wire  _sum_T_207 = tree_35_0_9 ^ tree_35_0_10; // @[Mul.scala 191:34]
  wire  ssum_2_17 = tree_35_0_9 ^ tree_35_0_10 ^ tree_35_0_11; // @[Mul.scala 191:42]
  wire  scout_2_17 = tree_35_0_9 & tree_35_0_10 | _sum_T_207 & tree_35_0_11; // @[Mul.scala 192:44]
  wire  _sum_T_209 = tree_35_0_12 ^ tree_35_0_13; // @[Mul.scala 191:34]
  wire  ssum_3_11 = tree_35_0_12 ^ tree_35_0_13 ^ tree_35_0_14; // @[Mul.scala 191:42]
  wire  scout_3_11 = tree_35_0_12 & tree_35_0_13 | _sum_T_209 & tree_35_0_14; // @[Mul.scala 192:44]
  wire  _sum_T_211 = tree_36_0 ^ tree_36_0_1; // @[Mul.scala 191:34]
  wire  sum_36 = tree_36_0 ^ tree_36_0_1 ^ tree_36_0_2; // @[Mul.scala 191:42]
  wire  cout_36 = tree_36_0 & tree_36_0_1 | _sum_T_211 & tree_36_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_213 = tree_36_0_3 ^ tree_36_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_28 = tree_36_0_3 ^ tree_36_0_4 ^ tree_36_0_5; // @[Mul.scala 191:42]
  wire  scout_0_28 = tree_36_0_3 & tree_36_0_4 | _sum_T_213 & tree_36_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_215 = tree_36_0_6 ^ tree_36_0_7; // @[Mul.scala 191:34]
  wire  ssum_1_24 = tree_36_0_6 ^ tree_36_0_7 ^ tree_36_0_8; // @[Mul.scala 191:42]
  wire  scout_1_24 = tree_36_0_6 & tree_36_0_7 | _sum_T_215 & tree_36_0_8; // @[Mul.scala 192:44]
  wire  _sum_T_217 = tree_36_0_9 ^ tree_36_0_10; // @[Mul.scala 191:34]
  wire  ssum_2_18 = tree_36_0_9 ^ tree_36_0_10 ^ tree_36_0_11; // @[Mul.scala 191:42]
  wire  scout_2_18 = tree_36_0_9 & tree_36_0_10 | _sum_T_217 & tree_36_0_11; // @[Mul.scala 192:44]
  wire  ssum_3_12 = tree_36_0_12 ^ tree_36_0_13; // @[Mul.scala 206:34]
  wire  scout_3_12 = tree_36_0_12 & tree_36_0_13; // @[Mul.scala 207:34]
  wire  _sum_T_220 = tree_37_0 ^ tree_37_0_1; // @[Mul.scala 191:34]
  wire  sum_37 = tree_37_0 ^ tree_37_0_1 ^ tree_37_0_2; // @[Mul.scala 191:42]
  wire  cout_37 = tree_37_0 & tree_37_0_1 | _sum_T_220 & tree_37_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_222 = tree_37_0_3 ^ tree_37_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_29 = tree_37_0_3 ^ tree_37_0_4 ^ tree_37_0_5; // @[Mul.scala 191:42]
  wire  scout_0_29 = tree_37_0_3 & tree_37_0_4 | _sum_T_222 & tree_37_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_224 = tree_37_0_6 ^ tree_37_0_7; // @[Mul.scala 191:34]
  wire  ssum_1_25 = tree_37_0_6 ^ tree_37_0_7 ^ tree_37_0_8; // @[Mul.scala 191:42]
  wire  scout_1_25 = tree_37_0_6 & tree_37_0_7 | _sum_T_224 & tree_37_0_8; // @[Mul.scala 192:44]
  wire  _sum_T_226 = tree_37_0_9 ^ tree_37_0_10; // @[Mul.scala 191:34]
  wire  ssum_2_19 = tree_37_0_9 ^ tree_37_0_10 ^ tree_37_0_11; // @[Mul.scala 191:42]
  wire  scout_2_19 = tree_37_0_9 & tree_37_0_10 | _sum_T_226 & tree_37_0_11; // @[Mul.scala 192:44]
  wire  ssum_3_13 = tree_37_0_12 ^ tree_37_0_13; // @[Mul.scala 206:34]
  wire  scout_3_13 = tree_37_0_12 & tree_37_0_13; // @[Mul.scala 207:34]
  wire  _sum_T_229 = tree_38_0 ^ tree_38_0_1; // @[Mul.scala 191:34]
  wire  sum_38 = tree_38_0 ^ tree_38_0_1 ^ tree_38_0_2; // @[Mul.scala 191:42]
  wire  cout_38 = tree_38_0 & tree_38_0_1 | _sum_T_229 & tree_38_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_231 = tree_38_0_3 ^ tree_38_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_30 = tree_38_0_3 ^ tree_38_0_4 ^ tree_38_0_5; // @[Mul.scala 191:42]
  wire  scout_0_30 = tree_38_0_3 & tree_38_0_4 | _sum_T_231 & tree_38_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_233 = tree_38_0_6 ^ tree_38_0_7; // @[Mul.scala 191:34]
  wire  ssum_1_26 = tree_38_0_6 ^ tree_38_0_7 ^ tree_38_0_8; // @[Mul.scala 191:42]
  wire  scout_1_26 = tree_38_0_6 & tree_38_0_7 | _sum_T_233 & tree_38_0_8; // @[Mul.scala 192:44]
  wire  ssum_2_20 = tree_38_0_9 ^ tree_38_0_10; // @[Mul.scala 206:34]
  wire  scout_2_20 = tree_38_0_9 & tree_38_0_10; // @[Mul.scala 207:34]
  wire  ssum_3_14 = tree_38_0_11 ^ tree_38_0_12; // @[Mul.scala 206:34]
  wire  scout_3_14 = tree_38_0_11 & tree_38_0_12; // @[Mul.scala 207:34]
  wire  _sum_T_237 = tree_39_0 ^ tree_39_0_1; // @[Mul.scala 191:34]
  wire  sum_39 = tree_39_0 ^ tree_39_0_1 ^ tree_39_0_2; // @[Mul.scala 191:42]
  wire  cout_39 = tree_39_0 & tree_39_0_1 | _sum_T_237 & tree_39_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_239 = tree_39_0_3 ^ tree_39_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_31 = tree_39_0_3 ^ tree_39_0_4 ^ tree_39_0_5; // @[Mul.scala 191:42]
  wire  scout_0_31 = tree_39_0_3 & tree_39_0_4 | _sum_T_239 & tree_39_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_241 = tree_39_0_6 ^ tree_39_0_7; // @[Mul.scala 191:34]
  wire  ssum_1_27 = tree_39_0_6 ^ tree_39_0_7 ^ tree_39_0_8; // @[Mul.scala 191:42]
  wire  scout_1_27 = tree_39_0_6 & tree_39_0_7 | _sum_T_241 & tree_39_0_8; // @[Mul.scala 192:44]
  wire  ssum_2_21 = tree_39_0_9 ^ tree_39_0_10; // @[Mul.scala 206:34]
  wire  scout_2_21 = tree_39_0_9 & tree_39_0_10; // @[Mul.scala 207:34]
  wire  ssum_3_15 = tree_39_0_11 ^ tree_39_0_12; // @[Mul.scala 206:34]
  wire  scout_3_15 = tree_39_0_11 & tree_39_0_12; // @[Mul.scala 207:34]
  wire  _sum_T_245 = tree_40_0 ^ tree_40_0_1; // @[Mul.scala 191:34]
  wire  sum_40 = tree_40_0 ^ tree_40_0_1 ^ tree_40_0_2; // @[Mul.scala 191:42]
  wire  cout_40 = tree_40_0 & tree_40_0_1 | _sum_T_245 & tree_40_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_247 = tree_40_0_3 ^ tree_40_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_32 = tree_40_0_3 ^ tree_40_0_4 ^ tree_40_0_5; // @[Mul.scala 191:42]
  wire  scout_0_32 = tree_40_0_3 & tree_40_0_4 | _sum_T_247 & tree_40_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_249 = tree_40_0_6 ^ tree_40_0_7; // @[Mul.scala 191:34]
  wire  ssum_1_28 = tree_40_0_6 ^ tree_40_0_7 ^ tree_40_0_8; // @[Mul.scala 191:42]
  wire  scout_1_28 = tree_40_0_6 & tree_40_0_7 | _sum_T_249 & tree_40_0_8; // @[Mul.scala 192:44]
  wire  _sum_T_251 = tree_40_0_9 ^ tree_40_0_10; // @[Mul.scala 191:34]
  wire  ssum_2_22 = tree_40_0_9 ^ tree_40_0_10 ^ tree_40_0_11; // @[Mul.scala 191:42]
  wire  scout_2_22 = tree_40_0_9 & tree_40_0_10 | _sum_T_251 & tree_40_0_11; // @[Mul.scala 192:44]
  wire  _sum_T_253 = tree_41_0 ^ tree_41_0_1; // @[Mul.scala 191:34]
  wire  sum_41 = tree_41_0 ^ tree_41_0_1 ^ tree_41_0_2; // @[Mul.scala 191:42]
  wire  cout_41 = tree_41_0 & tree_41_0_1 | _sum_T_253 & tree_41_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_255 = tree_41_0_3 ^ tree_41_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_33 = tree_41_0_3 ^ tree_41_0_4 ^ tree_41_0_5; // @[Mul.scala 191:42]
  wire  scout_0_33 = tree_41_0_3 & tree_41_0_4 | _sum_T_255 & tree_41_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_257 = tree_41_0_6 ^ tree_41_0_7; // @[Mul.scala 191:34]
  wire  ssum_1_29 = tree_41_0_6 ^ tree_41_0_7 ^ tree_41_0_8; // @[Mul.scala 191:42]
  wire  scout_1_29 = tree_41_0_6 & tree_41_0_7 | _sum_T_257 & tree_41_0_8; // @[Mul.scala 192:44]
  wire  _sum_T_259 = tree_41_0_9 ^ tree_41_0_10; // @[Mul.scala 191:34]
  wire  ssum_2_23 = tree_41_0_9 ^ tree_41_0_10 ^ tree_41_0_11; // @[Mul.scala 191:42]
  wire  scout_2_23 = tree_41_0_9 & tree_41_0_10 | _sum_T_259 & tree_41_0_11; // @[Mul.scala 192:44]
  wire  _sum_T_261 = tree_42_0 ^ tree_42_0_1; // @[Mul.scala 191:34]
  wire  sum_42 = tree_42_0 ^ tree_42_0_1 ^ tree_42_0_2; // @[Mul.scala 191:42]
  wire  cout_42 = tree_42_0 & tree_42_0_1 | _sum_T_261 & tree_42_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_263 = tree_42_0_3 ^ tree_42_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_34 = tree_42_0_3 ^ tree_42_0_4 ^ tree_42_0_5; // @[Mul.scala 191:42]
  wire  scout_0_34 = tree_42_0_3 & tree_42_0_4 | _sum_T_263 & tree_42_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_265 = tree_42_0_6 ^ tree_42_0_7; // @[Mul.scala 191:34]
  wire  ssum_1_30 = tree_42_0_6 ^ tree_42_0_7 ^ tree_42_0_8; // @[Mul.scala 191:42]
  wire  scout_1_30 = tree_42_0_6 & tree_42_0_7 | _sum_T_265 & tree_42_0_8; // @[Mul.scala 192:44]
  wire  ssum_2_24 = tree_42_0_9 ^ tree_42_0_10; // @[Mul.scala 206:34]
  wire  scout_2_24 = tree_42_0_9 & tree_42_0_10; // @[Mul.scala 207:34]
  wire  _sum_T_268 = tree_43_0 ^ tree_43_0_1; // @[Mul.scala 191:34]
  wire  sum_43 = tree_43_0 ^ tree_43_0_1 ^ tree_43_0_2; // @[Mul.scala 191:42]
  wire  cout_43 = tree_43_0 & tree_43_0_1 | _sum_T_268 & tree_43_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_270 = tree_43_0_3 ^ tree_43_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_35 = tree_43_0_3 ^ tree_43_0_4 ^ tree_43_0_5; // @[Mul.scala 191:42]
  wire  scout_0_35 = tree_43_0_3 & tree_43_0_4 | _sum_T_270 & tree_43_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_272 = tree_43_0_6 ^ tree_43_0_7; // @[Mul.scala 191:34]
  wire  ssum_1_31 = tree_43_0_6 ^ tree_43_0_7 ^ tree_43_0_8; // @[Mul.scala 191:42]
  wire  scout_1_31 = tree_43_0_6 & tree_43_0_7 | _sum_T_272 & tree_43_0_8; // @[Mul.scala 192:44]
  wire  ssum_2_25 = tree_43_0_9 ^ tree_43_0_10; // @[Mul.scala 206:34]
  wire  scout_2_25 = tree_43_0_9 & tree_43_0_10; // @[Mul.scala 207:34]
  wire  _sum_T_275 = tree_44_0 ^ tree_44_0_1; // @[Mul.scala 191:34]
  wire  sum_44 = tree_44_0 ^ tree_44_0_1 ^ tree_44_0_2; // @[Mul.scala 191:42]
  wire  cout_44 = tree_44_0 & tree_44_0_1 | _sum_T_275 & tree_44_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_277 = tree_44_0_3 ^ tree_44_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_36 = tree_44_0_3 ^ tree_44_0_4 ^ tree_44_0_5; // @[Mul.scala 191:42]
  wire  scout_0_36 = tree_44_0_3 & tree_44_0_4 | _sum_T_277 & tree_44_0_5; // @[Mul.scala 192:44]
  wire  ssum_1_32 = tree_44_0_6 ^ tree_44_0_7; // @[Mul.scala 206:34]
  wire  scout_1_32 = tree_44_0_6 & tree_44_0_7; // @[Mul.scala 207:34]
  wire  ssum_2_26 = tree_44_0_8 ^ tree_44_0_9; // @[Mul.scala 206:34]
  wire  scout_2_26 = tree_44_0_8 & tree_44_0_9; // @[Mul.scala 207:34]
  wire  _sum_T_281 = tree_45_0 ^ tree_45_0_1; // @[Mul.scala 191:34]
  wire  sum_45 = tree_45_0 ^ tree_45_0_1 ^ tree_45_0_2; // @[Mul.scala 191:42]
  wire  cout_45 = tree_45_0 & tree_45_0_1 | _sum_T_281 & tree_45_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_283 = tree_45_0_3 ^ tree_45_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_37 = tree_45_0_3 ^ tree_45_0_4 ^ tree_45_0_5; // @[Mul.scala 191:42]
  wire  scout_0_37 = tree_45_0_3 & tree_45_0_4 | _sum_T_283 & tree_45_0_5; // @[Mul.scala 192:44]
  wire  ssum_1_33 = tree_45_0_6 ^ tree_45_0_7; // @[Mul.scala 206:34]
  wire  scout_1_33 = tree_45_0_6 & tree_45_0_7; // @[Mul.scala 207:34]
  wire  ssum_2_27 = tree_45_0_8 ^ tree_45_0_9; // @[Mul.scala 206:34]
  wire  scout_2_27 = tree_45_0_8 & tree_45_0_9; // @[Mul.scala 207:34]
  wire  _sum_T_287 = tree_46_0 ^ tree_46_0_1; // @[Mul.scala 191:34]
  wire  sum_46 = tree_46_0 ^ tree_46_0_1 ^ tree_46_0_2; // @[Mul.scala 191:42]
  wire  cout_46 = tree_46_0 & tree_46_0_1 | _sum_T_287 & tree_46_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_289 = tree_46_0_3 ^ tree_46_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_38 = tree_46_0_3 ^ tree_46_0_4 ^ tree_46_0_5; // @[Mul.scala 191:42]
  wire  scout_0_38 = tree_46_0_3 & tree_46_0_4 | _sum_T_289 & tree_46_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_291 = tree_46_0_6 ^ tree_46_0_7; // @[Mul.scala 191:34]
  wire  ssum_1_34 = tree_46_0_6 ^ tree_46_0_7 ^ tree_46_0_8; // @[Mul.scala 191:42]
  wire  scout_1_34 = tree_46_0_6 & tree_46_0_7 | _sum_T_291 & tree_46_0_8; // @[Mul.scala 192:44]
  wire  _sum_T_293 = tree_47_0 ^ tree_47_0_1; // @[Mul.scala 191:34]
  wire  sum_47 = tree_47_0 ^ tree_47_0_1 ^ tree_47_0_2; // @[Mul.scala 191:42]
  wire  cout_47 = tree_47_0 & tree_47_0_1 | _sum_T_293 & tree_47_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_295 = tree_47_0_3 ^ tree_47_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_39 = tree_47_0_3 ^ tree_47_0_4 ^ tree_47_0_5; // @[Mul.scala 191:42]
  wire  scout_0_39 = tree_47_0_3 & tree_47_0_4 | _sum_T_295 & tree_47_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_297 = tree_47_0_6 ^ tree_47_0_7; // @[Mul.scala 191:34]
  wire  ssum_1_35 = tree_47_0_6 ^ tree_47_0_7 ^ tree_47_0_8; // @[Mul.scala 191:42]
  wire  scout_1_35 = tree_47_0_6 & tree_47_0_7 | _sum_T_297 & tree_47_0_8; // @[Mul.scala 192:44]
  wire  _sum_T_299 = tree_48_0 ^ tree_48_0_1; // @[Mul.scala 191:34]
  wire  sum_48 = tree_48_0 ^ tree_48_0_1 ^ tree_48_0_2; // @[Mul.scala 191:42]
  wire  cout_48 = tree_48_0 & tree_48_0_1 | _sum_T_299 & tree_48_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_301 = tree_48_0_3 ^ tree_48_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_40 = tree_48_0_3 ^ tree_48_0_4 ^ tree_48_0_5; // @[Mul.scala 191:42]
  wire  scout_0_40 = tree_48_0_3 & tree_48_0_4 | _sum_T_301 & tree_48_0_5; // @[Mul.scala 192:44]
  wire  ssum_1_36 = tree_48_0_6 ^ tree_48_0_7; // @[Mul.scala 206:34]
  wire  scout_1_36 = tree_48_0_6 & tree_48_0_7; // @[Mul.scala 207:34]
  wire  _sum_T_304 = tree_49_0 ^ tree_49_0_1; // @[Mul.scala 191:34]
  wire  sum_49 = tree_49_0 ^ tree_49_0_1 ^ tree_49_0_2; // @[Mul.scala 191:42]
  wire  cout_49 = tree_49_0 & tree_49_0_1 | _sum_T_304 & tree_49_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_306 = tree_49_0_3 ^ tree_49_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_41 = tree_49_0_3 ^ tree_49_0_4 ^ tree_49_0_5; // @[Mul.scala 191:42]
  wire  scout_0_41 = tree_49_0_3 & tree_49_0_4 | _sum_T_306 & tree_49_0_5; // @[Mul.scala 192:44]
  wire  ssum_1_37 = tree_49_0_6 ^ tree_49_0_7; // @[Mul.scala 206:34]
  wire  scout_1_37 = tree_49_0_6 & tree_49_0_7; // @[Mul.scala 207:34]
  wire  _sum_T_309 = tree_50_0 ^ tree_50_0_1; // @[Mul.scala 191:34]
  wire  sum_50 = tree_50_0 ^ tree_50_0_1 ^ tree_50_0_2; // @[Mul.scala 191:42]
  wire  cout_50 = tree_50_0 & tree_50_0_1 | _sum_T_309 & tree_50_0_2; // @[Mul.scala 192:44]
  wire  ssum_0_42 = tree_50_0_3 ^ tree_50_0_4; // @[Mul.scala 206:34]
  wire  scout_0_42 = tree_50_0_3 & tree_50_0_4; // @[Mul.scala 207:34]
  wire  ssum_1_38 = tree_50_0_5 ^ tree_50_0_6; // @[Mul.scala 206:34]
  wire  scout_1_38 = tree_50_0_5 & tree_50_0_6; // @[Mul.scala 207:34]
  wire  _sum_T_313 = tree_51_0 ^ tree_51_0_1; // @[Mul.scala 191:34]
  wire  sum_51 = tree_51_0 ^ tree_51_0_1 ^ tree_51_0_2; // @[Mul.scala 191:42]
  wire  cout_51 = tree_51_0 & tree_51_0_1 | _sum_T_313 & tree_51_0_2; // @[Mul.scala 192:44]
  wire  ssum_0_43 = tree_51_0_3 ^ tree_51_0_4; // @[Mul.scala 206:34]
  wire  scout_0_43 = tree_51_0_3 & tree_51_0_4; // @[Mul.scala 207:34]
  wire  ssum_1_39 = tree_51_0_5 ^ tree_51_0_6; // @[Mul.scala 206:34]
  wire  scout_1_39 = tree_51_0_5 & tree_51_0_6; // @[Mul.scala 207:34]
  wire  _sum_T_317 = tree_52_0 ^ tree_52_0_1; // @[Mul.scala 191:34]
  wire  sum_52 = tree_52_0 ^ tree_52_0_1 ^ tree_52_0_2; // @[Mul.scala 191:42]
  wire  cout_52 = tree_52_0 & tree_52_0_1 | _sum_T_317 & tree_52_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_319 = tree_52_0_3 ^ tree_52_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_44 = tree_52_0_3 ^ tree_52_0_4 ^ tree_52_0_5; // @[Mul.scala 191:42]
  wire  scout_0_44 = tree_52_0_3 & tree_52_0_4 | _sum_T_319 & tree_52_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_321 = tree_53_0 ^ tree_53_0_1; // @[Mul.scala 191:34]
  wire  sum_53 = tree_53_0 ^ tree_53_0_1 ^ tree_53_0_2; // @[Mul.scala 191:42]
  wire  cout_53 = tree_53_0 & tree_53_0_1 | _sum_T_321 & tree_53_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_323 = tree_53_0_3 ^ tree_53_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_45 = tree_53_0_3 ^ tree_53_0_4 ^ tree_53_0_5; // @[Mul.scala 191:42]
  wire  scout_0_45 = tree_53_0_3 & tree_53_0_4 | _sum_T_323 & tree_53_0_5; // @[Mul.scala 192:44]
  wire  _sum_T_325 = tree_54_0 ^ tree_54_0_1; // @[Mul.scala 191:34]
  wire  sum_54 = tree_54_0 ^ tree_54_0_1 ^ tree_54_0_2; // @[Mul.scala 191:42]
  wire  cout_54 = tree_54_0 & tree_54_0_1 | _sum_T_325 & tree_54_0_2; // @[Mul.scala 192:44]
  wire  ssum_0_46 = tree_54_0_3 ^ tree_54_0_4; // @[Mul.scala 206:34]
  wire  scout_0_46 = tree_54_0_3 & tree_54_0_4; // @[Mul.scala 207:34]
  wire  _sum_T_328 = tree_55_0 ^ tree_55_0_1; // @[Mul.scala 191:34]
  wire  sum_55 = tree_55_0 ^ tree_55_0_1 ^ tree_55_0_2; // @[Mul.scala 191:42]
  wire  cout_55 = tree_55_0 & tree_55_0_1 | _sum_T_328 & tree_55_0_2; // @[Mul.scala 192:44]
  wire  ssum_0_47 = tree_55_0_3 ^ tree_55_0_4; // @[Mul.scala 206:34]
  wire  scout_0_47 = tree_55_0_3 & tree_55_0_4; // @[Mul.scala 207:34]
  wire  sum_56 = tree_56_0 ^ tree_56_0_1; // @[Mul.scala 206:34]
  wire  cout_56 = tree_56_0 & tree_56_0_1; // @[Mul.scala 207:34]
  wire  sum_57 = tree_56_0_2 ^ tree_56_0_3; // @[Mul.scala 206:34]
  wire  cout_57 = tree_56_0_2 & tree_56_0_3; // @[Mul.scala 207:34]
  wire  sum_58 = tree_57_0 ^ tree_57_0_1; // @[Mul.scala 206:34]
  wire  cout_58 = tree_57_0 & tree_57_0_1; // @[Mul.scala 207:34]
  wire  sum_59 = tree_57_0_2 ^ tree_57_0_3; // @[Mul.scala 206:34]
  wire  cout_59 = tree_57_0_2 & tree_57_0_3; // @[Mul.scala 207:34]
  wire  _sum_T_335 = tree_58_0 ^ tree_58_0_1; // @[Mul.scala 191:34]
  wire  sum_60 = tree_58_0 ^ tree_58_0_1 ^ tree_58_0_2; // @[Mul.scala 191:42]
  wire  cout_60 = tree_58_0 & tree_58_0_1 | _sum_T_335 & tree_58_0_2; // @[Mul.scala 192:44]
  wire  _sum_T_337 = tree_59_0 ^ tree_59_0_1; // @[Mul.scala 191:34]
  wire  sum_61 = tree_59_0 ^ tree_59_0_1 ^ tree_59_0_2; // @[Mul.scala 191:42]
  wire  cout_61 = tree_59_0 & tree_59_0_1 | _sum_T_337 & tree_59_0_2; // @[Mul.scala 192:44]
  wire  sum_62 = tree_60_0 ^ tree_60_0_1; // @[Mul.scala 206:34]
  wire  cout_62 = tree_60_0 & tree_60_0_1; // @[Mul.scala 207:34]
  wire  sum_63 = tree_61_0 ^ tree_61_0_1; // @[Mul.scala 206:34]
  wire  cout_63 = tree_61_0 & tree_61_0_1; // @[Mul.scala 207:34]
  wire  sum_66 = sum_1 ^ cout; // @[Mul.scala 206:34]
  wire  cout_66 = sum_1 & cout; // @[Mul.scala 207:34]
  wire  sum_67 = sum_2 ^ cout_1; // @[Mul.scala 206:34]
  wire  cout_67 = sum_2 & cout_1; // @[Mul.scala 207:34]
  wire  sum_68 = sum_3 ^ cout_2; // @[Mul.scala 206:34]
  wire  cout_68 = sum_3 & cout_2; // @[Mul.scala 207:34]
  wire  _sum_T_346 = sum_4 ^ sum_5; // @[Mul.scala 191:34]
  wire  sum_69 = sum_4 ^ sum_5 ^ cout_3; // @[Mul.scala 191:42]
  wire  cout_69 = sum_4 & sum_5 | _sum_T_346 & cout_3; // @[Mul.scala 192:44]
  wire  sum_70 = sum_6 ^ sum_7; // @[Mul.scala 206:34]
  wire  cout_70 = sum_6 & sum_7; // @[Mul.scala 207:34]
  wire  sum_71 = cout_4 ^ cout_5; // @[Mul.scala 206:34]
  wire  cout_71 = cout_4 & cout_5; // @[Mul.scala 207:34]
  wire  sum_72 = sum_8 ^ ssum_0; // @[Mul.scala 206:34]
  wire  cout_72 = sum_8 & ssum_0; // @[Mul.scala 207:34]
  wire  sum_73 = cout_6 ^ cout_7; // @[Mul.scala 206:34]
  wire  cout_73 = cout_6 & cout_7; // @[Mul.scala 207:34]
  wire  sum_74 = sum_9 ^ ssum_0_1; // @[Mul.scala 206:34]
  wire  cout_74 = sum_9 & ssum_0_1; // @[Mul.scala 207:34]
  wire  sum_75 = cout_8 ^ scout_0; // @[Mul.scala 206:34]
  wire  cout_75 = cout_8 & scout_0; // @[Mul.scala 207:34]
  wire  sum_76 = sum_10 ^ ssum_0_2; // @[Mul.scala 206:34]
  wire  cout_76 = sum_10 & ssum_0_2; // @[Mul.scala 207:34]
  wire  sum_77 = cout_9 ^ scout_0_1; // @[Mul.scala 206:34]
  wire  cout_77 = cout_9 & scout_0_1; // @[Mul.scala 207:34]
  wire  sum_78 = sum_11 ^ ssum_0_3; // @[Mul.scala 206:34]
  wire  cout_78 = sum_11 & ssum_0_3; // @[Mul.scala 207:34]
  wire  sum_79 = cout_10 ^ scout_0_2; // @[Mul.scala 206:34]
  wire  cout_79 = cout_10 & scout_0_2; // @[Mul.scala 207:34]
  wire  _sum_T_358 = sum_12 ^ ssum_0_4; // @[Mul.scala 191:34]
  wire  sum_80 = sum_12 ^ ssum_0_4 ^ ssum_1; // @[Mul.scala 191:42]
  wire  cout_80 = sum_12 & ssum_0_4 | _sum_T_358 & ssum_1; // @[Mul.scala 192:44]
  wire  ssum_0_48 = cout_11 ^ scout_0_3; // @[Mul.scala 206:34]
  wire  scout_0_48 = cout_11 & scout_0_3; // @[Mul.scala 207:34]
  wire  _sum_T_361 = sum_13 ^ ssum_0_5; // @[Mul.scala 191:34]
  wire  sum_81 = sum_13 ^ ssum_0_5 ^ ssum_1_1; // @[Mul.scala 191:42]
  wire  cout_81 = sum_13 & ssum_0_5 | _sum_T_361 & ssum_1_1; // @[Mul.scala 192:44]
  wire  _sum_T_363 = cout_12 ^ scout_0_4; // @[Mul.scala 191:34]
  wire  ssum_0_49 = cout_12 ^ scout_0_4 ^ scout_1; // @[Mul.scala 191:42]
  wire  scout_0_49 = cout_12 & scout_0_4 | _sum_T_363 & scout_1; // @[Mul.scala 192:44]
  wire  _sum_T_365 = sum_14 ^ ssum_0_6; // @[Mul.scala 191:34]
  wire  sum_82 = sum_14 ^ ssum_0_6 ^ ssum_1_2; // @[Mul.scala 191:42]
  wire  cout_82 = sum_14 & ssum_0_6 | _sum_T_365 & ssum_1_2; // @[Mul.scala 192:44]
  wire  _sum_T_367 = cout_13 ^ scout_0_5; // @[Mul.scala 191:34]
  wire  ssum_0_50 = cout_13 ^ scout_0_5 ^ scout_1_1; // @[Mul.scala 191:42]
  wire  scout_0_50 = cout_13 & scout_0_5 | _sum_T_367 & scout_1_1; // @[Mul.scala 192:44]
  wire  _sum_T_369 = sum_15 ^ ssum_0_7; // @[Mul.scala 191:34]
  wire  sum_83 = sum_15 ^ ssum_0_7 ^ ssum_1_3; // @[Mul.scala 191:42]
  wire  cout_83 = sum_15 & ssum_0_7 | _sum_T_369 & ssum_1_3; // @[Mul.scala 192:44]
  wire  _sum_T_371 = cout_14 ^ scout_0_6; // @[Mul.scala 191:34]
  wire  ssum_0_51 = cout_14 ^ scout_0_6 ^ scout_1_2; // @[Mul.scala 191:42]
  wire  scout_0_51 = cout_14 & scout_0_6 | _sum_T_371 & scout_1_2; // @[Mul.scala 192:44]
  wire  _sum_T_373 = sum_16 ^ ssum_0_8; // @[Mul.scala 191:34]
  wire  sum_84 = sum_16 ^ ssum_0_8 ^ ssum_1_4; // @[Mul.scala 191:42]
  wire  cout_84 = sum_16 & ssum_0_8 | _sum_T_373 & ssum_1_4; // @[Mul.scala 192:44]
  wire  _sum_T_375 = cout_15 ^ scout_0_7; // @[Mul.scala 191:34]
  wire  ssum_0_52 = cout_15 ^ scout_0_7 ^ scout_1_3; // @[Mul.scala 191:42]
  wire  scout_0_52 = cout_15 & scout_0_7 | _sum_T_375 & scout_1_3; // @[Mul.scala 192:44]
  wire  _sum_T_377 = sum_17 ^ ssum_0_9; // @[Mul.scala 191:34]
  wire  sum_85 = sum_17 ^ ssum_0_9 ^ ssum_1_5; // @[Mul.scala 191:42]
  wire  cout_85 = sum_17 & ssum_0_9 | _sum_T_377 & ssum_1_5; // @[Mul.scala 192:44]
  wire  _sum_T_379 = cout_16 ^ scout_0_8; // @[Mul.scala 191:34]
  wire  ssum_0_53 = cout_16 ^ scout_0_8 ^ scout_1_4; // @[Mul.scala 191:42]
  wire  scout_0_53 = cout_16 & scout_0_8 | _sum_T_379 & scout_1_4; // @[Mul.scala 192:44]
  wire  _sum_T_381 = sum_18 ^ ssum_0_10; // @[Mul.scala 191:34]
  wire  sum_86 = sum_18 ^ ssum_0_10 ^ ssum_1_6; // @[Mul.scala 191:42]
  wire  cout_86 = sum_18 & ssum_0_10 | _sum_T_381 & ssum_1_6; // @[Mul.scala 192:44]
  wire  ssum_0_54 = ssum_2 ^ cout_17; // @[Mul.scala 206:34]
  wire  scout_0_54 = ssum_2 & cout_17; // @[Mul.scala 207:34]
  wire  ssum_1_40 = scout_0_9 ^ scout_1_5; // @[Mul.scala 206:34]
  wire  scout_1_40 = scout_0_9 & scout_1_5; // @[Mul.scala 207:34]
  wire  _sum_T_385 = sum_19 ^ ssum_0_11; // @[Mul.scala 191:34]
  wire  sum_87 = sum_19 ^ ssum_0_11 ^ ssum_1_7; // @[Mul.scala 191:42]
  wire  cout_87 = sum_19 & ssum_0_11 | _sum_T_385 & ssum_1_7; // @[Mul.scala 192:44]
  wire  _sum_T_387 = ssum_2_1 ^ cout_18; // @[Mul.scala 191:34]
  wire  ssum_0_55 = ssum_2_1 ^ cout_18 ^ scout_0_10; // @[Mul.scala 191:42]
  wire  scout_0_55 = ssum_2_1 & cout_18 | _sum_T_387 & scout_0_10; // @[Mul.scala 192:44]
  wire  ssum_1_41 = scout_1_6 ^ scout_2; // @[Mul.scala 206:34]
  wire  scout_1_41 = scout_1_6 & scout_2; // @[Mul.scala 207:34]
  wire  _sum_T_390 = sum_20 ^ ssum_0_12; // @[Mul.scala 191:34]
  wire  sum_88 = sum_20 ^ ssum_0_12 ^ ssum_1_8; // @[Mul.scala 191:42]
  wire  cout_88 = sum_20 & ssum_0_12 | _sum_T_390 & ssum_1_8; // @[Mul.scala 192:44]
  wire  _sum_T_392 = ssum_2_2 ^ cout_19; // @[Mul.scala 191:34]
  wire  ssum_0_56 = ssum_2_2 ^ cout_19 ^ scout_0_11; // @[Mul.scala 191:42]
  wire  scout_0_56 = ssum_2_2 & cout_19 | _sum_T_392 & scout_0_11; // @[Mul.scala 192:44]
  wire  ssum_1_42 = scout_1_7 ^ scout_2_1; // @[Mul.scala 206:34]
  wire  scout_1_42 = scout_1_7 & scout_2_1; // @[Mul.scala 207:34]
  wire  _sum_T_395 = sum_21 ^ ssum_0_13; // @[Mul.scala 191:34]
  wire  sum_89 = sum_21 ^ ssum_0_13 ^ ssum_1_9; // @[Mul.scala 191:42]
  wire  cout_89 = sum_21 & ssum_0_13 | _sum_T_395 & ssum_1_9; // @[Mul.scala 192:44]
  wire  _sum_T_397 = ssum_2_3 ^ cout_20; // @[Mul.scala 191:34]
  wire  ssum_0_57 = ssum_2_3 ^ cout_20 ^ scout_0_12; // @[Mul.scala 191:42]
  wire  scout_0_57 = ssum_2_3 & cout_20 | _sum_T_397 & scout_0_12; // @[Mul.scala 192:44]
  wire  ssum_1_43 = scout_1_8 ^ scout_2_2; // @[Mul.scala 206:34]
  wire  scout_1_43 = scout_1_8 & scout_2_2; // @[Mul.scala 207:34]
  wire  _sum_T_400 = sum_22 ^ ssum_0_14; // @[Mul.scala 191:34]
  wire  sum_90 = sum_22 ^ ssum_0_14 ^ ssum_1_10; // @[Mul.scala 191:42]
  wire  cout_90 = sum_22 & ssum_0_14 | _sum_T_400 & ssum_1_10; // @[Mul.scala 192:44]
  wire  _sum_T_402 = ssum_2_4 ^ cout_21; // @[Mul.scala 191:34]
  wire  ssum_0_58 = ssum_2_4 ^ cout_21 ^ scout_0_13; // @[Mul.scala 191:42]
  wire  scout_0_58 = ssum_2_4 & cout_21 | _sum_T_402 & scout_0_13; // @[Mul.scala 192:44]
  wire  ssum_1_44 = scout_1_9 ^ scout_2_3; // @[Mul.scala 206:34]
  wire  scout_1_44 = scout_1_9 & scout_2_3; // @[Mul.scala 207:34]
  wire  _sum_T_405 = sum_23 ^ ssum_0_15; // @[Mul.scala 191:34]
  wire  sum_91 = sum_23 ^ ssum_0_15 ^ ssum_1_11; // @[Mul.scala 191:42]
  wire  cout_91 = sum_23 & ssum_0_15 | _sum_T_405 & ssum_1_11; // @[Mul.scala 192:44]
  wire  _sum_T_407 = ssum_2_5 ^ cout_22; // @[Mul.scala 191:34]
  wire  ssum_0_59 = ssum_2_5 ^ cout_22 ^ scout_0_14; // @[Mul.scala 191:42]
  wire  scout_0_59 = ssum_2_5 & cout_22 | _sum_T_407 & scout_0_14; // @[Mul.scala 192:44]
  wire  ssum_1_45 = scout_1_10 ^ scout_2_4; // @[Mul.scala 206:34]
  wire  scout_1_45 = scout_1_10 & scout_2_4; // @[Mul.scala 207:34]
  wire  _sum_T_410 = sum_24 ^ ssum_0_16; // @[Mul.scala 191:34]
  wire  sum_92 = sum_24 ^ ssum_0_16 ^ ssum_1_12; // @[Mul.scala 191:42]
  wire  cout_92 = sum_24 & ssum_0_16 | _sum_T_410 & ssum_1_12; // @[Mul.scala 192:44]
  wire  _sum_T_412 = ssum_2_6 ^ ssum_3; // @[Mul.scala 191:34]
  wire  ssum_0_60 = ssum_2_6 ^ ssum_3 ^ cout_23; // @[Mul.scala 191:42]
  wire  scout_0_60 = ssum_2_6 & ssum_3 | _sum_T_412 & cout_23; // @[Mul.scala 192:44]
  wire  _sum_T_414 = scout_0_15 ^ scout_1_11; // @[Mul.scala 191:34]
  wire  ssum_1_46 = scout_0_15 ^ scout_1_11 ^ scout_2_5; // @[Mul.scala 191:42]
  wire  scout_1_46 = scout_0_15 & scout_1_11 | _sum_T_414 & scout_2_5; // @[Mul.scala 192:44]
  wire  _sum_T_416 = sum_25 ^ ssum_0_17; // @[Mul.scala 191:34]
  wire  sum_93 = sum_25 ^ ssum_0_17 ^ ssum_1_13; // @[Mul.scala 191:42]
  wire  cout_93 = sum_25 & ssum_0_17 | _sum_T_416 & ssum_1_13; // @[Mul.scala 192:44]
  wire  _sum_T_418 = ssum_2_7 ^ ssum_3_1; // @[Mul.scala 191:34]
  wire  ssum_0_61 = ssum_2_7 ^ ssum_3_1 ^ cout_24; // @[Mul.scala 191:42]
  wire  scout_0_61 = ssum_2_7 & ssum_3_1 | _sum_T_418 & cout_24; // @[Mul.scala 192:44]
  wire  ssum_1_47 = scout_0_16 ^ scout_1_12; // @[Mul.scala 206:34]
  wire  scout_1_47 = scout_0_16 & scout_1_12; // @[Mul.scala 207:34]
  wire  ssum_2_28 = scout_2_6 ^ scout_3; // @[Mul.scala 206:34]
  wire  scout_2_28 = scout_2_6 & scout_3; // @[Mul.scala 207:34]
  wire  _sum_T_422 = sum_26 ^ ssum_0_18; // @[Mul.scala 191:34]
  wire  sum_94 = sum_26 ^ ssum_0_18 ^ ssum_1_14; // @[Mul.scala 191:42]
  wire  cout_94 = sum_26 & ssum_0_18 | _sum_T_422 & ssum_1_14; // @[Mul.scala 192:44]
  wire  _sum_T_424 = ssum_2_8 ^ ssum_3_2; // @[Mul.scala 191:34]
  wire  ssum_0_62 = ssum_2_8 ^ ssum_3_2 ^ cout_25; // @[Mul.scala 191:42]
  wire  scout_0_62 = ssum_2_8 & ssum_3_2 | _sum_T_424 & cout_25; // @[Mul.scala 192:44]
  wire  ssum_1_48 = scout_0_17 ^ scout_1_13; // @[Mul.scala 206:34]
  wire  scout_1_48 = scout_0_17 & scout_1_13; // @[Mul.scala 207:34]
  wire  ssum_2_29 = scout_2_7 ^ scout_3_1; // @[Mul.scala 206:34]
  wire  scout_2_29 = scout_2_7 & scout_3_1; // @[Mul.scala 207:34]
  wire  _sum_T_428 = sum_27 ^ ssum_0_19; // @[Mul.scala 191:34]
  wire  sum_95 = sum_27 ^ ssum_0_19 ^ ssum_1_15; // @[Mul.scala 191:42]
  wire  cout_95 = sum_27 & ssum_0_19 | _sum_T_428 & ssum_1_15; // @[Mul.scala 192:44]
  wire  _sum_T_430 = ssum_2_9 ^ ssum_3_3; // @[Mul.scala 191:34]
  wire  ssum_0_63 = ssum_2_9 ^ ssum_3_3 ^ cout_26; // @[Mul.scala 191:42]
  wire  scout_0_63 = ssum_2_9 & ssum_3_3 | _sum_T_430 & cout_26; // @[Mul.scala 192:44]
  wire  ssum_1_49 = scout_0_18 ^ scout_1_14; // @[Mul.scala 206:34]
  wire  scout_1_49 = scout_0_18 & scout_1_14; // @[Mul.scala 207:34]
  wire  ssum_2_30 = scout_2_8 ^ scout_3_2; // @[Mul.scala 206:34]
  wire  scout_2_30 = scout_2_8 & scout_3_2; // @[Mul.scala 207:34]
  wire  _sum_T_434 = sum_28 ^ ssum_0_20; // @[Mul.scala 191:34]
  wire  sum_96 = sum_28 ^ ssum_0_20 ^ ssum_1_16; // @[Mul.scala 191:42]
  wire  cout_96 = sum_28 & ssum_0_20 | _sum_T_434 & ssum_1_16; // @[Mul.scala 192:44]
  wire  _sum_T_436 = ssum_2_10 ^ ssum_3_4; // @[Mul.scala 191:34]
  wire  ssum_0_64 = ssum_2_10 ^ ssum_3_4 ^ cout_27; // @[Mul.scala 191:42]
  wire  scout_0_64 = ssum_2_10 & ssum_3_4 | _sum_T_436 & cout_27; // @[Mul.scala 192:44]
  wire  ssum_1_50 = scout_0_19 ^ scout_1_15; // @[Mul.scala 206:34]
  wire  scout_1_50 = scout_0_19 & scout_1_15; // @[Mul.scala 207:34]
  wire  ssum_2_31 = scout_2_9 ^ scout_3_3; // @[Mul.scala 206:34]
  wire  scout_2_31 = scout_2_9 & scout_3_3; // @[Mul.scala 207:34]
  wire  _sum_T_440 = sum_29 ^ ssum_0_21; // @[Mul.scala 191:34]
  wire  sum_97 = sum_29 ^ ssum_0_21 ^ ssum_1_17; // @[Mul.scala 191:42]
  wire  cout_97 = sum_29 & ssum_0_21 | _sum_T_440 & ssum_1_17; // @[Mul.scala 192:44]
  wire  _sum_T_442 = ssum_2_11 ^ ssum_3_5; // @[Mul.scala 191:34]
  wire  ssum_0_65 = ssum_2_11 ^ ssum_3_5 ^ cout_28; // @[Mul.scala 191:42]
  wire  scout_0_65 = ssum_2_11 & ssum_3_5 | _sum_T_442 & cout_28; // @[Mul.scala 192:44]
  wire  ssum_1_51 = scout_0_20 ^ scout_1_16; // @[Mul.scala 206:34]
  wire  scout_1_51 = scout_0_20 & scout_1_16; // @[Mul.scala 207:34]
  wire  ssum_2_32 = scout_2_10 ^ scout_3_4; // @[Mul.scala 206:34]
  wire  scout_2_32 = scout_2_10 & scout_3_4; // @[Mul.scala 207:34]
  wire  _sum_T_446 = sum_30 ^ ssum_0_22; // @[Mul.scala 191:34]
  wire  sum_98 = sum_30 ^ ssum_0_22 ^ ssum_1_18; // @[Mul.scala 191:42]
  wire  cout_98 = sum_30 & ssum_0_22 | _sum_T_446 & ssum_1_18; // @[Mul.scala 192:44]
  wire  _sum_T_448 = ssum_2_12 ^ ssum_3_6; // @[Mul.scala 191:34]
  wire  ssum_0_66 = ssum_2_12 ^ ssum_3_6 ^ ssum_4; // @[Mul.scala 191:42]
  wire  scout_0_66 = ssum_2_12 & ssum_3_6 | _sum_T_448 & ssum_4; // @[Mul.scala 192:44]
  wire  _sum_T_450 = cout_29 ^ scout_0_21; // @[Mul.scala 191:34]
  wire  ssum_1_52 = cout_29 ^ scout_0_21 ^ scout_1_17; // @[Mul.scala 191:42]
  wire  scout_1_52 = cout_29 & scout_0_21 | _sum_T_450 & scout_1_17; // @[Mul.scala 192:44]
  wire  ssum_2_33 = scout_2_11 ^ scout_3_5; // @[Mul.scala 206:34]
  wire  scout_2_33 = scout_2_11 & scout_3_5; // @[Mul.scala 207:34]
  wire  _sum_T_453 = sum_31 ^ ssum_0_23; // @[Mul.scala 191:34]
  wire  sum_99 = sum_31 ^ ssum_0_23 ^ ssum_1_19; // @[Mul.scala 191:42]
  wire  cout_99 = sum_31 & ssum_0_23 | _sum_T_453 & ssum_1_19; // @[Mul.scala 192:44]
  wire  _sum_T_455 = ssum_2_13 ^ ssum_3_7; // @[Mul.scala 191:34]
  wire  ssum_0_67 = ssum_2_13 ^ ssum_3_7 ^ ssum_4_1; // @[Mul.scala 191:42]
  wire  scout_0_67 = ssum_2_13 & ssum_3_7 | _sum_T_455 & ssum_4_1; // @[Mul.scala 192:44]
  wire  _sum_T_457 = cout_30 ^ scout_0_22; // @[Mul.scala 191:34]
  wire  ssum_1_53 = cout_30 ^ scout_0_22 ^ scout_1_18; // @[Mul.scala 191:42]
  wire  scout_1_53 = cout_30 & scout_0_22 | _sum_T_457 & scout_1_18; // @[Mul.scala 192:44]
  wire  _sum_T_459 = scout_2_12 ^ scout_3_6; // @[Mul.scala 191:34]
  wire  ssum_2_34 = scout_2_12 ^ scout_3_6 ^ scout_4; // @[Mul.scala 191:42]
  wire  scout_2_34 = scout_2_12 & scout_3_6 | _sum_T_459 & scout_4; // @[Mul.scala 192:44]
  wire  _sum_T_461 = sum_32 ^ ssum_0_24; // @[Mul.scala 191:34]
  wire  sum_100 = sum_32 ^ ssum_0_24 ^ ssum_1_20; // @[Mul.scala 191:42]
  wire  cout_100 = sum_32 & ssum_0_24 | _sum_T_461 & ssum_1_20; // @[Mul.scala 192:44]
  wire  _sum_T_463 = ssum_2_14 ^ ssum_3_8; // @[Mul.scala 191:34]
  wire  ssum_0_68 = ssum_2_14 ^ ssum_3_8 ^ ssum_4_2; // @[Mul.scala 191:42]
  wire  scout_0_68 = ssum_2_14 & ssum_3_8 | _sum_T_463 & ssum_4_2; // @[Mul.scala 192:44]
  wire  _sum_T_465 = cout_31 ^ scout_0_23; // @[Mul.scala 191:34]
  wire  ssum_1_54 = cout_31 ^ scout_0_23 ^ scout_1_19; // @[Mul.scala 191:42]
  wire  scout_1_54 = cout_31 & scout_0_23 | _sum_T_465 & scout_1_19; // @[Mul.scala 192:44]
  wire  _sum_T_467 = scout_2_13 ^ scout_3_7; // @[Mul.scala 191:34]
  wire  ssum_2_35 = scout_2_13 ^ scout_3_7 ^ scout_4_1; // @[Mul.scala 191:42]
  wire  scout_2_35 = scout_2_13 & scout_3_7 | _sum_T_467 & scout_4_1; // @[Mul.scala 192:44]
  wire  _sum_T_469 = sum_33 ^ ssum_0_25; // @[Mul.scala 191:34]
  wire  sum_101 = sum_33 ^ ssum_0_25 ^ ssum_1_21; // @[Mul.scala 191:42]
  wire  cout_101 = sum_33 & ssum_0_25 | _sum_T_469 & ssum_1_21; // @[Mul.scala 192:44]
  wire  _sum_T_471 = ssum_2_15 ^ ssum_3_9; // @[Mul.scala 191:34]
  wire  ssum_0_69 = ssum_2_15 ^ ssum_3_9 ^ ssum_4_3; // @[Mul.scala 191:42]
  wire  scout_0_69 = ssum_2_15 & ssum_3_9 | _sum_T_471 & ssum_4_3; // @[Mul.scala 192:44]
  wire  _sum_T_473 = cout_32 ^ scout_0_24; // @[Mul.scala 191:34]
  wire  ssum_1_55 = cout_32 ^ scout_0_24 ^ scout_1_20; // @[Mul.scala 191:42]
  wire  scout_1_55 = cout_32 & scout_0_24 | _sum_T_473 & scout_1_20; // @[Mul.scala 192:44]
  wire  _sum_T_475 = scout_2_14 ^ scout_3_8; // @[Mul.scala 191:34]
  wire  ssum_2_36 = scout_2_14 ^ scout_3_8 ^ tree_32_0_15; // @[Mul.scala 191:42]
  wire  scout_2_36 = scout_2_14 & scout_3_8 | _sum_T_475 & tree_32_0_15; // @[Mul.scala 192:44]
  wire  _sum_T_477 = sum_34 ^ ssum_0_26; // @[Mul.scala 191:34]
  wire  sum_102 = sum_34 ^ ssum_0_26 ^ ssum_1_22; // @[Mul.scala 191:42]
  wire  cout_102 = sum_34 & ssum_0_26 | _sum_T_477 & ssum_1_22; // @[Mul.scala 192:44]
  wire  _sum_T_479 = ssum_2_16 ^ ssum_3_10; // @[Mul.scala 191:34]
  wire  ssum_0_70 = ssum_2_16 ^ ssum_3_10 ^ cout_33; // @[Mul.scala 191:42]
  wire  scout_0_70 = ssum_2_16 & ssum_3_10 | _sum_T_479 & cout_33; // @[Mul.scala 192:44]
  wire  _sum_T_481 = scout_0_25 ^ scout_1_21; // @[Mul.scala 191:34]
  wire  ssum_1_56 = scout_0_25 ^ scout_1_21 ^ scout_2_15; // @[Mul.scala 191:42]
  wire  scout_1_56 = scout_0_25 & scout_1_21 | _sum_T_481 & scout_2_15; // @[Mul.scala 192:44]
  wire  ssum_2_37 = scout_3_9 ^ scout_4_3; // @[Mul.scala 206:34]
  wire  scout_2_37 = scout_3_9 & scout_4_3; // @[Mul.scala 207:34]
  wire  _sum_T_484 = sum_35 ^ ssum_0_27; // @[Mul.scala 191:34]
  wire  sum_103 = sum_35 ^ ssum_0_27 ^ ssum_1_23; // @[Mul.scala 191:42]
  wire  cout_103 = sum_35 & ssum_0_27 | _sum_T_484 & ssum_1_23; // @[Mul.scala 192:44]
  wire  _sum_T_486 = ssum_2_17 ^ ssum_3_11; // @[Mul.scala 191:34]
  wire  ssum_0_71 = ssum_2_17 ^ ssum_3_11 ^ cout_34; // @[Mul.scala 191:42]
  wire  scout_0_71 = ssum_2_17 & ssum_3_11 | _sum_T_486 & cout_34; // @[Mul.scala 192:44]
  wire  ssum_1_57 = scout_0_26 ^ scout_1_22; // @[Mul.scala 206:34]
  wire  scout_1_57 = scout_0_26 & scout_1_22; // @[Mul.scala 207:34]
  wire  ssum_2_38 = scout_2_16 ^ scout_3_10; // @[Mul.scala 206:34]
  wire  scout_2_38 = scout_2_16 & scout_3_10; // @[Mul.scala 207:34]
  wire  _sum_T_490 = sum_36 ^ ssum_0_28; // @[Mul.scala 191:34]
  wire  sum_104 = sum_36 ^ ssum_0_28 ^ ssum_1_24; // @[Mul.scala 191:42]
  wire  cout_104 = sum_36 & ssum_0_28 | _sum_T_490 & ssum_1_24; // @[Mul.scala 192:44]
  wire  _sum_T_492 = ssum_2_18 ^ ssum_3_12; // @[Mul.scala 191:34]
  wire  ssum_0_72 = ssum_2_18 ^ ssum_3_12 ^ cout_35; // @[Mul.scala 191:42]
  wire  scout_0_72 = ssum_2_18 & ssum_3_12 | _sum_T_492 & cout_35; // @[Mul.scala 192:44]
  wire  ssum_1_58 = scout_0_27 ^ scout_1_23; // @[Mul.scala 206:34]
  wire  scout_1_58 = scout_0_27 & scout_1_23; // @[Mul.scala 207:34]
  wire  ssum_2_39 = scout_2_17 ^ scout_3_11; // @[Mul.scala 206:34]
  wire  scout_2_39 = scout_2_17 & scout_3_11; // @[Mul.scala 207:34]
  wire  _sum_T_496 = sum_37 ^ ssum_0_29; // @[Mul.scala 191:34]
  wire  sum_105 = sum_37 ^ ssum_0_29 ^ ssum_1_25; // @[Mul.scala 191:42]
  wire  cout_105 = sum_37 & ssum_0_29 | _sum_T_496 & ssum_1_25; // @[Mul.scala 192:44]
  wire  _sum_T_498 = ssum_2_19 ^ ssum_3_13; // @[Mul.scala 191:34]
  wire  ssum_0_73 = ssum_2_19 ^ ssum_3_13 ^ cout_36; // @[Mul.scala 191:42]
  wire  scout_0_73 = ssum_2_19 & ssum_3_13 | _sum_T_498 & cout_36; // @[Mul.scala 192:44]
  wire  ssum_1_59 = scout_0_28 ^ scout_1_24; // @[Mul.scala 206:34]
  wire  scout_1_59 = scout_0_28 & scout_1_24; // @[Mul.scala 207:34]
  wire  ssum_2_40 = scout_2_18 ^ scout_3_12; // @[Mul.scala 206:34]
  wire  scout_2_40 = scout_2_18 & scout_3_12; // @[Mul.scala 207:34]
  wire  _sum_T_502 = sum_38 ^ ssum_0_30; // @[Mul.scala 191:34]
  wire  sum_106 = sum_38 ^ ssum_0_30 ^ ssum_1_26; // @[Mul.scala 191:42]
  wire  cout_106 = sum_38 & ssum_0_30 | _sum_T_502 & ssum_1_26; // @[Mul.scala 192:44]
  wire  _sum_T_504 = ssum_2_20 ^ ssum_3_14; // @[Mul.scala 191:34]
  wire  ssum_0_74 = ssum_2_20 ^ ssum_3_14 ^ cout_37; // @[Mul.scala 191:42]
  wire  scout_0_74 = ssum_2_20 & ssum_3_14 | _sum_T_504 & cout_37; // @[Mul.scala 192:44]
  wire  ssum_1_60 = scout_0_29 ^ scout_1_25; // @[Mul.scala 206:34]
  wire  scout_1_60 = scout_0_29 & scout_1_25; // @[Mul.scala 207:34]
  wire  ssum_2_41 = scout_2_19 ^ scout_3_13; // @[Mul.scala 206:34]
  wire  scout_2_41 = scout_2_19 & scout_3_13; // @[Mul.scala 207:34]
  wire  _sum_T_508 = sum_39 ^ ssum_0_31; // @[Mul.scala 191:34]
  wire  sum_107 = sum_39 ^ ssum_0_31 ^ ssum_1_27; // @[Mul.scala 191:42]
  wire  cout_107 = sum_39 & ssum_0_31 | _sum_T_508 & ssum_1_27; // @[Mul.scala 192:44]
  wire  _sum_T_510 = ssum_2_21 ^ ssum_3_15; // @[Mul.scala 191:34]
  wire  ssum_0_75 = ssum_2_21 ^ ssum_3_15 ^ cout_38; // @[Mul.scala 191:42]
  wire  scout_0_75 = ssum_2_21 & ssum_3_15 | _sum_T_510 & cout_38; // @[Mul.scala 192:44]
  wire  ssum_1_61 = scout_0_30 ^ scout_1_26; // @[Mul.scala 206:34]
  wire  scout_1_61 = scout_0_30 & scout_1_26; // @[Mul.scala 207:34]
  wire  ssum_2_42 = scout_2_20 ^ scout_3_14; // @[Mul.scala 206:34]
  wire  scout_2_42 = scout_2_20 & scout_3_14; // @[Mul.scala 207:34]
  wire  _sum_T_514 = sum_40 ^ ssum_0_32; // @[Mul.scala 191:34]
  wire  sum_108 = sum_40 ^ ssum_0_32 ^ ssum_1_28; // @[Mul.scala 191:42]
  wire  cout_108 = sum_40 & ssum_0_32 | _sum_T_514 & ssum_1_28; // @[Mul.scala 192:44]
  wire  _sum_T_516 = ssum_2_22 ^ cout_39; // @[Mul.scala 191:34]
  wire  ssum_0_76 = ssum_2_22 ^ cout_39 ^ scout_0_31; // @[Mul.scala 191:42]
  wire  scout_0_76 = ssum_2_22 & cout_39 | _sum_T_516 & scout_0_31; // @[Mul.scala 192:44]
  wire  _sum_T_518 = scout_1_27 ^ scout_2_21; // @[Mul.scala 191:34]
  wire  ssum_1_62 = scout_1_27 ^ scout_2_21 ^ scout_3_15; // @[Mul.scala 191:42]
  wire  scout_1_62 = scout_1_27 & scout_2_21 | _sum_T_518 & scout_3_15; // @[Mul.scala 192:44]
  wire  _sum_T_520 = sum_41 ^ ssum_0_33; // @[Mul.scala 191:34]
  wire  sum_109 = sum_41 ^ ssum_0_33 ^ ssum_1_29; // @[Mul.scala 191:42]
  wire  cout_109 = sum_41 & ssum_0_33 | _sum_T_520 & ssum_1_29; // @[Mul.scala 192:44]
  wire  _sum_T_522 = ssum_2_23 ^ cout_40; // @[Mul.scala 191:34]
  wire  ssum_0_77 = ssum_2_23 ^ cout_40 ^ scout_0_32; // @[Mul.scala 191:42]
  wire  scout_0_77 = ssum_2_23 & cout_40 | _sum_T_522 & scout_0_32; // @[Mul.scala 192:44]
  wire  ssum_1_63 = scout_1_28 ^ scout_2_22; // @[Mul.scala 206:34]
  wire  scout_1_63 = scout_1_28 & scout_2_22; // @[Mul.scala 207:34]
  wire  _sum_T_525 = sum_42 ^ ssum_0_34; // @[Mul.scala 191:34]
  wire  sum_110 = sum_42 ^ ssum_0_34 ^ ssum_1_30; // @[Mul.scala 191:42]
  wire  cout_110 = sum_42 & ssum_0_34 | _sum_T_525 & ssum_1_30; // @[Mul.scala 192:44]
  wire  _sum_T_527 = ssum_2_24 ^ cout_41; // @[Mul.scala 191:34]
  wire  ssum_0_78 = ssum_2_24 ^ cout_41 ^ scout_0_33; // @[Mul.scala 191:42]
  wire  scout_0_78 = ssum_2_24 & cout_41 | _sum_T_527 & scout_0_33; // @[Mul.scala 192:44]
  wire  ssum_1_64 = scout_1_29 ^ scout_2_23; // @[Mul.scala 206:34]
  wire  scout_1_64 = scout_1_29 & scout_2_23; // @[Mul.scala 207:34]
  wire  _sum_T_530 = sum_43 ^ ssum_0_35; // @[Mul.scala 191:34]
  wire  sum_111 = sum_43 ^ ssum_0_35 ^ ssum_1_31; // @[Mul.scala 191:42]
  wire  cout_111 = sum_43 & ssum_0_35 | _sum_T_530 & ssum_1_31; // @[Mul.scala 192:44]
  wire  _sum_T_532 = ssum_2_25 ^ cout_42; // @[Mul.scala 191:34]
  wire  ssum_0_79 = ssum_2_25 ^ cout_42 ^ scout_0_34; // @[Mul.scala 191:42]
  wire  scout_0_79 = ssum_2_25 & cout_42 | _sum_T_532 & scout_0_34; // @[Mul.scala 192:44]
  wire  ssum_1_65 = scout_1_30 ^ scout_2_24; // @[Mul.scala 206:34]
  wire  scout_1_65 = scout_1_30 & scout_2_24; // @[Mul.scala 207:34]
  wire  _sum_T_535 = sum_44 ^ ssum_0_36; // @[Mul.scala 191:34]
  wire  sum_112 = sum_44 ^ ssum_0_36 ^ ssum_1_32; // @[Mul.scala 191:42]
  wire  cout_112 = sum_44 & ssum_0_36 | _sum_T_535 & ssum_1_32; // @[Mul.scala 192:44]
  wire  _sum_T_537 = ssum_2_26 ^ cout_43; // @[Mul.scala 191:34]
  wire  ssum_0_80 = ssum_2_26 ^ cout_43 ^ scout_0_35; // @[Mul.scala 191:42]
  wire  scout_0_80 = ssum_2_26 & cout_43 | _sum_T_537 & scout_0_35; // @[Mul.scala 192:44]
  wire  ssum_1_66 = scout_1_31 ^ scout_2_25; // @[Mul.scala 206:34]
  wire  scout_1_66 = scout_1_31 & scout_2_25; // @[Mul.scala 207:34]
  wire  _sum_T_540 = sum_45 ^ ssum_0_37; // @[Mul.scala 191:34]
  wire  sum_113 = sum_45 ^ ssum_0_37 ^ ssum_1_33; // @[Mul.scala 191:42]
  wire  cout_113 = sum_45 & ssum_0_37 | _sum_T_540 & ssum_1_33; // @[Mul.scala 192:44]
  wire  _sum_T_542 = ssum_2_27 ^ cout_44; // @[Mul.scala 191:34]
  wire  ssum_0_81 = ssum_2_27 ^ cout_44 ^ scout_0_36; // @[Mul.scala 191:42]
  wire  scout_0_81 = ssum_2_27 & cout_44 | _sum_T_542 & scout_0_36; // @[Mul.scala 192:44]
  wire  ssum_1_67 = scout_1_32 ^ scout_2_26; // @[Mul.scala 206:34]
  wire  scout_1_67 = scout_1_32 & scout_2_26; // @[Mul.scala 207:34]
  wire  _sum_T_545 = sum_46 ^ ssum_0_38; // @[Mul.scala 191:34]
  wire  sum_114 = sum_46 ^ ssum_0_38 ^ ssum_1_34; // @[Mul.scala 191:42]
  wire  cout_114 = sum_46 & ssum_0_38 | _sum_T_545 & ssum_1_34; // @[Mul.scala 192:44]
  wire  ssum_0_82 = cout_45 ^ scout_0_37; // @[Mul.scala 206:34]
  wire  scout_0_82 = cout_45 & scout_0_37; // @[Mul.scala 207:34]
  wire  ssum_1_68 = scout_1_33 ^ scout_2_27; // @[Mul.scala 206:34]
  wire  scout_1_68 = scout_1_33 & scout_2_27; // @[Mul.scala 207:34]
  wire  _sum_T_549 = sum_47 ^ ssum_0_39; // @[Mul.scala 191:34]
  wire  sum_115 = sum_47 ^ ssum_0_39 ^ ssum_1_35; // @[Mul.scala 191:42]
  wire  cout_115 = sum_47 & ssum_0_39 | _sum_T_549 & ssum_1_35; // @[Mul.scala 192:44]
  wire  _sum_T_551 = cout_46 ^ scout_0_38; // @[Mul.scala 191:34]
  wire  ssum_0_83 = cout_46 ^ scout_0_38 ^ scout_1_34; // @[Mul.scala 191:42]
  wire  scout_0_83 = cout_46 & scout_0_38 | _sum_T_551 & scout_1_34; // @[Mul.scala 192:44]
  wire  _sum_T_553 = sum_48 ^ ssum_0_40; // @[Mul.scala 191:34]
  wire  sum_116 = sum_48 ^ ssum_0_40 ^ ssum_1_36; // @[Mul.scala 191:42]
  wire  cout_116 = sum_48 & ssum_0_40 | _sum_T_553 & ssum_1_36; // @[Mul.scala 192:44]
  wire  _sum_T_555 = cout_47 ^ scout_0_39; // @[Mul.scala 191:34]
  wire  ssum_0_84 = cout_47 ^ scout_0_39 ^ scout_1_35; // @[Mul.scala 191:42]
  wire  scout_0_84 = cout_47 & scout_0_39 | _sum_T_555 & scout_1_35; // @[Mul.scala 192:44]
  wire  _sum_T_557 = sum_49 ^ ssum_0_41; // @[Mul.scala 191:34]
  wire  sum_117 = sum_49 ^ ssum_0_41 ^ ssum_1_37; // @[Mul.scala 191:42]
  wire  cout_117 = sum_49 & ssum_0_41 | _sum_T_557 & ssum_1_37; // @[Mul.scala 192:44]
  wire  _sum_T_559 = cout_48 ^ scout_0_40; // @[Mul.scala 191:34]
  wire  ssum_0_85 = cout_48 ^ scout_0_40 ^ scout_1_36; // @[Mul.scala 191:42]
  wire  scout_0_85 = cout_48 & scout_0_40 | _sum_T_559 & scout_1_36; // @[Mul.scala 192:44]
  wire  _sum_T_561 = sum_50 ^ ssum_0_42; // @[Mul.scala 191:34]
  wire  sum_118 = sum_50 ^ ssum_0_42 ^ ssum_1_38; // @[Mul.scala 191:42]
  wire  cout_118 = sum_50 & ssum_0_42 | _sum_T_561 & ssum_1_38; // @[Mul.scala 192:44]
  wire  _sum_T_563 = cout_49 ^ scout_0_41; // @[Mul.scala 191:34]
  wire  ssum_0_86 = cout_49 ^ scout_0_41 ^ scout_1_37; // @[Mul.scala 191:42]
  wire  scout_0_86 = cout_49 & scout_0_41 | _sum_T_563 & scout_1_37; // @[Mul.scala 192:44]
  wire  _sum_T_565 = sum_51 ^ ssum_0_43; // @[Mul.scala 191:34]
  wire  sum_119 = sum_51 ^ ssum_0_43 ^ ssum_1_39; // @[Mul.scala 191:42]
  wire  cout_119 = sum_51 & ssum_0_43 | _sum_T_565 & ssum_1_39; // @[Mul.scala 192:44]
  wire  _sum_T_567 = cout_50 ^ scout_0_42; // @[Mul.scala 191:34]
  wire  ssum_0_87 = cout_50 ^ scout_0_42 ^ scout_1_38; // @[Mul.scala 191:42]
  wire  scout_0_87 = cout_50 & scout_0_42 | _sum_T_567 & scout_1_38; // @[Mul.scala 192:44]
  wire  _sum_T_569 = sum_52 ^ ssum_0_44; // @[Mul.scala 191:34]
  wire  sum_120 = sum_52 ^ ssum_0_44 ^ cout_51; // @[Mul.scala 191:42]
  wire  cout_120 = sum_52 & ssum_0_44 | _sum_T_569 & cout_51; // @[Mul.scala 192:44]
  wire  ssum_0_88 = scout_0_43 ^ scout_1_39; // @[Mul.scala 206:34]
  wire  scout_0_88 = scout_0_43 & scout_1_39; // @[Mul.scala 207:34]
  wire  sum_121 = sum_53 ^ ssum_0_45; // @[Mul.scala 206:34]
  wire  cout_121 = sum_53 & ssum_0_45; // @[Mul.scala 207:34]
  wire  sum_122 = cout_52 ^ scout_0_44; // @[Mul.scala 206:34]
  wire  cout_122 = cout_52 & scout_0_44; // @[Mul.scala 207:34]
  wire  sum_123 = sum_54 ^ ssum_0_46; // @[Mul.scala 206:34]
  wire  cout_123 = sum_54 & ssum_0_46; // @[Mul.scala 207:34]
  wire  sum_124 = cout_53 ^ scout_0_45; // @[Mul.scala 206:34]
  wire  cout_124 = cout_53 & scout_0_45; // @[Mul.scala 207:34]
  wire  sum_125 = sum_55 ^ ssum_0_47; // @[Mul.scala 206:34]
  wire  cout_125 = sum_55 & ssum_0_47; // @[Mul.scala 207:34]
  wire  sum_126 = cout_54 ^ scout_0_46; // @[Mul.scala 206:34]
  wire  cout_126 = cout_54 & scout_0_46; // @[Mul.scala 207:34]
  wire  sum_127 = sum_56 ^ sum_57; // @[Mul.scala 206:34]
  wire  cout_127 = sum_56 & sum_57; // @[Mul.scala 207:34]
  wire  sum_128 = cout_55 ^ scout_0_47; // @[Mul.scala 206:34]
  wire  cout_128 = cout_55 & scout_0_47; // @[Mul.scala 207:34]
  wire  sum_129 = sum_58 ^ sum_59; // @[Mul.scala 206:34]
  wire  cout_129 = sum_58 & sum_59; // @[Mul.scala 207:34]
  wire  sum_130 = cout_56 ^ cout_57; // @[Mul.scala 206:34]
  wire  cout_130 = cout_56 & cout_57; // @[Mul.scala 207:34]
  wire  _sum_T_582 = sum_60 ^ cout_58; // @[Mul.scala 191:34]
  wire  sum_131 = sum_60 ^ cout_58 ^ cout_59; // @[Mul.scala 191:42]
  wire  cout_131 = sum_60 & cout_58 | _sum_T_582 & cout_59; // @[Mul.scala 192:44]
  wire  sum_132 = sum_61 ^ cout_60; // @[Mul.scala 206:34]
  wire  cout_132 = sum_61 & cout_60; // @[Mul.scala 207:34]
  wire  sum_133 = sum_62 ^ cout_61; // @[Mul.scala 206:34]
  wire  cout_133 = sum_62 & cout_61; // @[Mul.scala 207:34]
  wire  sum_134 = sum_63 ^ cout_62; // @[Mul.scala 206:34]
  wire  cout_134 = sum_63 & cout_62; // @[Mul.scala 207:34]
  wire  sum_135 = tree_62_0 ^ cout_63; // @[Mul.scala 206:34]
  wire  cout_135 = tree_62_0 & cout_63; // @[Mul.scala 207:34]
  wire  sum_140 = sum_67 ^ cout_66; // @[Mul.scala 206:34]
  wire  cout_140 = sum_67 & cout_66; // @[Mul.scala 207:34]
  wire  sum_141 = sum_68 ^ cout_67; // @[Mul.scala 206:34]
  wire  cout_141 = sum_68 & cout_67; // @[Mul.scala 207:34]
  wire  sum_142 = sum_69 ^ cout_68; // @[Mul.scala 206:34]
  wire  cout_142 = sum_69 & cout_68; // @[Mul.scala 207:34]
  wire  _sum_T_595 = sum_70 ^ sum_71; // @[Mul.scala 191:34]
  wire  sum_143 = sum_70 ^ sum_71 ^ cout_69; // @[Mul.scala 191:42]
  wire  cout_143 = sum_70 & sum_71 | _sum_T_595 & cout_69; // @[Mul.scala 192:44]
  wire  sum_144 = sum_72 ^ sum_73; // @[Mul.scala 206:34]
  wire  cout_144 = sum_72 & sum_73; // @[Mul.scala 207:34]
  wire  sum_145 = cout_70 ^ cout_71; // @[Mul.scala 206:34]
  wire  cout_145 = cout_70 & cout_71; // @[Mul.scala 207:34]
  wire  sum_146 = sum_74 ^ sum_75; // @[Mul.scala 206:34]
  wire  cout_146 = sum_74 & sum_75; // @[Mul.scala 207:34]
  wire  sum_147 = cout_72 ^ cout_73; // @[Mul.scala 206:34]
  wire  cout_147 = cout_72 & cout_73; // @[Mul.scala 207:34]
  wire  sum_148 = sum_76 ^ sum_77; // @[Mul.scala 206:34]
  wire  cout_148 = sum_76 & sum_77; // @[Mul.scala 207:34]
  wire  sum_149 = cout_74 ^ cout_75; // @[Mul.scala 206:34]
  wire  cout_149 = cout_74 & cout_75; // @[Mul.scala 207:34]
  wire  sum_150 = sum_78 ^ sum_79; // @[Mul.scala 206:34]
  wire  cout_150 = sum_78 & sum_79; // @[Mul.scala 207:34]
  wire  sum_151 = cout_76 ^ cout_77; // @[Mul.scala 206:34]
  wire  cout_151 = cout_76 & cout_77; // @[Mul.scala 207:34]
  wire  sum_152 = sum_80 ^ ssum_0_48; // @[Mul.scala 206:34]
  wire  cout_152 = sum_80 & ssum_0_48; // @[Mul.scala 207:34]
  wire  sum_153 = cout_78 ^ cout_79; // @[Mul.scala 206:34]
  wire  cout_153 = cout_78 & cout_79; // @[Mul.scala 207:34]
  wire  sum_154 = sum_81 ^ ssum_0_49; // @[Mul.scala 206:34]
  wire  cout_154 = sum_81 & ssum_0_49; // @[Mul.scala 207:34]
  wire  sum_155 = cout_80 ^ scout_0_48; // @[Mul.scala 206:34]
  wire  cout_155 = cout_80 & scout_0_48; // @[Mul.scala 207:34]
  wire  sum_156 = sum_82 ^ ssum_0_50; // @[Mul.scala 206:34]
  wire  cout_156 = sum_82 & ssum_0_50; // @[Mul.scala 207:34]
  wire  sum_157 = cout_81 ^ scout_0_49; // @[Mul.scala 206:34]
  wire  cout_157 = cout_81 & scout_0_49; // @[Mul.scala 207:34]
  wire  sum_158 = sum_83 ^ ssum_0_51; // @[Mul.scala 206:34]
  wire  cout_158 = sum_83 & ssum_0_51; // @[Mul.scala 207:34]
  wire  sum_159 = cout_82 ^ scout_0_50; // @[Mul.scala 206:34]
  wire  cout_159 = cout_82 & scout_0_50; // @[Mul.scala 207:34]
  wire  sum_160 = sum_84 ^ ssum_0_52; // @[Mul.scala 206:34]
  wire  cout_160 = sum_84 & ssum_0_52; // @[Mul.scala 207:34]
  wire  sum_161 = cout_83 ^ scout_0_51; // @[Mul.scala 206:34]
  wire  cout_161 = cout_83 & scout_0_51; // @[Mul.scala 207:34]
  wire  sum_162 = sum_85 ^ ssum_0_53; // @[Mul.scala 206:34]
  wire  cout_162 = sum_85 & ssum_0_53; // @[Mul.scala 207:34]
  wire  sum_163 = cout_84 ^ scout_0_52; // @[Mul.scala 206:34]
  wire  cout_163 = cout_84 & scout_0_52; // @[Mul.scala 207:34]
  wire  _sum_T_617 = sum_86 ^ ssum_0_54; // @[Mul.scala 191:34]
  wire  sum_164 = sum_86 ^ ssum_0_54 ^ ssum_1_40; // @[Mul.scala 191:42]
  wire  cout_164 = sum_86 & ssum_0_54 | _sum_T_617 & ssum_1_40; // @[Mul.scala 192:44]
  wire  ssum_0_89 = cout_85 ^ scout_0_53; // @[Mul.scala 206:34]
  wire  scout_0_89 = cout_85 & scout_0_53; // @[Mul.scala 207:34]
  wire  _sum_T_620 = sum_87 ^ ssum_0_55; // @[Mul.scala 191:34]
  wire  sum_165 = sum_87 ^ ssum_0_55 ^ ssum_1_41; // @[Mul.scala 191:42]
  wire  cout_165 = sum_87 & ssum_0_55 | _sum_T_620 & ssum_1_41; // @[Mul.scala 192:44]
  wire  _sum_T_622 = cout_86 ^ scout_0_54; // @[Mul.scala 191:34]
  wire  ssum_0_90 = cout_86 ^ scout_0_54 ^ scout_1_40; // @[Mul.scala 191:42]
  wire  scout_0_90 = cout_86 & scout_0_54 | _sum_T_622 & scout_1_40; // @[Mul.scala 192:44]
  wire  _sum_T_624 = sum_88 ^ ssum_0_56; // @[Mul.scala 191:34]
  wire  sum_166 = sum_88 ^ ssum_0_56 ^ ssum_1_42; // @[Mul.scala 191:42]
  wire  cout_166 = sum_88 & ssum_0_56 | _sum_T_624 & ssum_1_42; // @[Mul.scala 192:44]
  wire  _sum_T_626 = cout_87 ^ scout_0_55; // @[Mul.scala 191:34]
  wire  ssum_0_91 = cout_87 ^ scout_0_55 ^ scout_1_41; // @[Mul.scala 191:42]
  wire  scout_0_91 = cout_87 & scout_0_55 | _sum_T_626 & scout_1_41; // @[Mul.scala 192:44]
  wire  _sum_T_628 = sum_89 ^ ssum_0_57; // @[Mul.scala 191:34]
  wire  sum_167 = sum_89 ^ ssum_0_57 ^ ssum_1_43; // @[Mul.scala 191:42]
  wire  cout_167 = sum_89 & ssum_0_57 | _sum_T_628 & ssum_1_43; // @[Mul.scala 192:44]
  wire  _sum_T_630 = cout_88 ^ scout_0_56; // @[Mul.scala 191:34]
  wire  ssum_0_92 = cout_88 ^ scout_0_56 ^ scout_1_42; // @[Mul.scala 191:42]
  wire  scout_0_92 = cout_88 & scout_0_56 | _sum_T_630 & scout_1_42; // @[Mul.scala 192:44]
  wire  _sum_T_632 = sum_90 ^ ssum_0_58; // @[Mul.scala 191:34]
  wire  sum_168 = sum_90 ^ ssum_0_58 ^ ssum_1_44; // @[Mul.scala 191:42]
  wire  cout_168 = sum_90 & ssum_0_58 | _sum_T_632 & ssum_1_44; // @[Mul.scala 192:44]
  wire  _sum_T_634 = cout_89 ^ scout_0_57; // @[Mul.scala 191:34]
  wire  ssum_0_93 = cout_89 ^ scout_0_57 ^ scout_1_43; // @[Mul.scala 191:42]
  wire  scout_0_93 = cout_89 & scout_0_57 | _sum_T_634 & scout_1_43; // @[Mul.scala 192:44]
  wire  _sum_T_636 = sum_91 ^ ssum_0_59; // @[Mul.scala 191:34]
  wire  sum_169 = sum_91 ^ ssum_0_59 ^ ssum_1_45; // @[Mul.scala 191:42]
  wire  cout_169 = sum_91 & ssum_0_59 | _sum_T_636 & ssum_1_45; // @[Mul.scala 192:44]
  wire  _sum_T_638 = cout_90 ^ scout_0_58; // @[Mul.scala 191:34]
  wire  ssum_0_94 = cout_90 ^ scout_0_58 ^ scout_1_44; // @[Mul.scala 191:42]
  wire  scout_0_94 = cout_90 & scout_0_58 | _sum_T_638 & scout_1_44; // @[Mul.scala 192:44]
  wire  _sum_T_640 = sum_92 ^ ssum_0_60; // @[Mul.scala 191:34]
  wire  sum_170 = sum_92 ^ ssum_0_60 ^ ssum_1_46; // @[Mul.scala 191:42]
  wire  cout_170 = sum_92 & ssum_0_60 | _sum_T_640 & ssum_1_46; // @[Mul.scala 192:44]
  wire  _sum_T_642 = cout_91 ^ scout_0_59; // @[Mul.scala 191:34]
  wire  ssum_0_95 = cout_91 ^ scout_0_59 ^ scout_1_45; // @[Mul.scala 191:42]
  wire  scout_0_95 = cout_91 & scout_0_59 | _sum_T_642 & scout_1_45; // @[Mul.scala 192:44]
  wire  _sum_T_644 = sum_93 ^ ssum_0_61; // @[Mul.scala 191:34]
  wire  sum_171 = sum_93 ^ ssum_0_61 ^ ssum_1_47; // @[Mul.scala 191:42]
  wire  cout_171 = sum_93 & ssum_0_61 | _sum_T_644 & ssum_1_47; // @[Mul.scala 192:44]
  wire  ssum_0_96 = ssum_2_28 ^ cout_92; // @[Mul.scala 206:34]
  wire  scout_0_96 = ssum_2_28 & cout_92; // @[Mul.scala 207:34]
  wire  ssum_1_69 = scout_0_60 ^ scout_1_46; // @[Mul.scala 206:34]
  wire  scout_1_69 = scout_0_60 & scout_1_46; // @[Mul.scala 207:34]
  wire  _sum_T_648 = sum_94 ^ ssum_0_62; // @[Mul.scala 191:34]
  wire  sum_172 = sum_94 ^ ssum_0_62 ^ ssum_1_48; // @[Mul.scala 191:42]
  wire  cout_172 = sum_94 & ssum_0_62 | _sum_T_648 & ssum_1_48; // @[Mul.scala 192:44]
  wire  _sum_T_650 = ssum_2_29 ^ cout_93; // @[Mul.scala 191:34]
  wire  ssum_0_97 = ssum_2_29 ^ cout_93 ^ scout_0_61; // @[Mul.scala 191:42]
  wire  scout_0_97 = ssum_2_29 & cout_93 | _sum_T_650 & scout_0_61; // @[Mul.scala 192:44]
  wire  ssum_1_70 = scout_1_47 ^ scout_2_28; // @[Mul.scala 206:34]
  wire  scout_1_70 = scout_1_47 & scout_2_28; // @[Mul.scala 207:34]
  wire  _sum_T_653 = sum_95 ^ ssum_0_63; // @[Mul.scala 191:34]
  wire  sum_173 = sum_95 ^ ssum_0_63 ^ ssum_1_49; // @[Mul.scala 191:42]
  wire  cout_173 = sum_95 & ssum_0_63 | _sum_T_653 & ssum_1_49; // @[Mul.scala 192:44]
  wire  _sum_T_655 = ssum_2_30 ^ cout_94; // @[Mul.scala 191:34]
  wire  ssum_0_98 = ssum_2_30 ^ cout_94 ^ scout_0_62; // @[Mul.scala 191:42]
  wire  scout_0_98 = ssum_2_30 & cout_94 | _sum_T_655 & scout_0_62; // @[Mul.scala 192:44]
  wire  ssum_1_71 = scout_1_48 ^ scout_2_29; // @[Mul.scala 206:34]
  wire  scout_1_71 = scout_1_48 & scout_2_29; // @[Mul.scala 207:34]
  wire  _sum_T_658 = sum_96 ^ ssum_0_64; // @[Mul.scala 191:34]
  wire  sum_174 = sum_96 ^ ssum_0_64 ^ ssum_1_50; // @[Mul.scala 191:42]
  wire  cout_174 = sum_96 & ssum_0_64 | _sum_T_658 & ssum_1_50; // @[Mul.scala 192:44]
  wire  _sum_T_660 = ssum_2_31 ^ cout_95; // @[Mul.scala 191:34]
  wire  ssum_0_99 = ssum_2_31 ^ cout_95 ^ scout_0_63; // @[Mul.scala 191:42]
  wire  scout_0_99 = ssum_2_31 & cout_95 | _sum_T_660 & scout_0_63; // @[Mul.scala 192:44]
  wire  ssum_1_72 = scout_1_49 ^ scout_2_30; // @[Mul.scala 206:34]
  wire  scout_1_72 = scout_1_49 & scout_2_30; // @[Mul.scala 207:34]
  wire  _sum_T_663 = sum_97 ^ ssum_0_65; // @[Mul.scala 191:34]
  wire  sum_175 = sum_97 ^ ssum_0_65 ^ ssum_1_51; // @[Mul.scala 191:42]
  wire  cout_175 = sum_97 & ssum_0_65 | _sum_T_663 & ssum_1_51; // @[Mul.scala 192:44]
  wire  _sum_T_665 = ssum_2_32 ^ cout_96; // @[Mul.scala 191:34]
  wire  ssum_0_100 = ssum_2_32 ^ cout_96 ^ scout_0_64; // @[Mul.scala 191:42]
  wire  scout_0_100 = ssum_2_32 & cout_96 | _sum_T_665 & scout_0_64; // @[Mul.scala 192:44]
  wire  ssum_1_73 = scout_1_50 ^ scout_2_31; // @[Mul.scala 206:34]
  wire  scout_1_73 = scout_1_50 & scout_2_31; // @[Mul.scala 207:34]
  wire  _sum_T_668 = sum_98 ^ ssum_0_66; // @[Mul.scala 191:34]
  wire  sum_176 = sum_98 ^ ssum_0_66 ^ ssum_1_52; // @[Mul.scala 191:42]
  wire  cout_176 = sum_98 & ssum_0_66 | _sum_T_668 & ssum_1_52; // @[Mul.scala 192:44]
  wire  _sum_T_670 = ssum_2_33 ^ cout_97; // @[Mul.scala 191:34]
  wire  ssum_0_101 = ssum_2_33 ^ cout_97 ^ scout_0_65; // @[Mul.scala 191:42]
  wire  scout_0_101 = ssum_2_33 & cout_97 | _sum_T_670 & scout_0_65; // @[Mul.scala 192:44]
  wire  ssum_1_74 = scout_1_51 ^ scout_2_32; // @[Mul.scala 206:34]
  wire  scout_1_74 = scout_1_51 & scout_2_32; // @[Mul.scala 207:34]
  wire  _sum_T_673 = sum_99 ^ ssum_0_67; // @[Mul.scala 191:34]
  wire  sum_177 = sum_99 ^ ssum_0_67 ^ ssum_1_53; // @[Mul.scala 191:42]
  wire  cout_177 = sum_99 & ssum_0_67 | _sum_T_673 & ssum_1_53; // @[Mul.scala 192:44]
  wire  _sum_T_675 = ssum_2_34 ^ cout_98; // @[Mul.scala 191:34]
  wire  ssum_0_102 = ssum_2_34 ^ cout_98 ^ scout_0_66; // @[Mul.scala 191:42]
  wire  scout_0_102 = ssum_2_34 & cout_98 | _sum_T_675 & scout_0_66; // @[Mul.scala 192:44]
  wire  ssum_1_75 = scout_1_52 ^ scout_2_33; // @[Mul.scala 206:34]
  wire  scout_1_75 = scout_1_52 & scout_2_33; // @[Mul.scala 207:34]
  wire  _sum_T_678 = sum_100 ^ ssum_0_68; // @[Mul.scala 191:34]
  wire  sum_178 = sum_100 ^ ssum_0_68 ^ ssum_1_54; // @[Mul.scala 191:42]
  wire  cout_178 = sum_100 & ssum_0_68 | _sum_T_678 & ssum_1_54; // @[Mul.scala 192:44]
  wire  _sum_T_680 = ssum_2_35 ^ cout_99; // @[Mul.scala 191:34]
  wire  ssum_0_103 = ssum_2_35 ^ cout_99 ^ scout_0_67; // @[Mul.scala 191:42]
  wire  scout_0_103 = ssum_2_35 & cout_99 | _sum_T_680 & scout_0_67; // @[Mul.scala 192:44]
  wire  ssum_1_76 = scout_1_53 ^ scout_2_34; // @[Mul.scala 206:34]
  wire  scout_1_76 = scout_1_53 & scout_2_34; // @[Mul.scala 207:34]
  wire  _sum_T_683 = sum_101 ^ ssum_0_69; // @[Mul.scala 191:34]
  wire  sum_179 = sum_101 ^ ssum_0_69 ^ ssum_1_55; // @[Mul.scala 191:42]
  wire  cout_179 = sum_101 & ssum_0_69 | _sum_T_683 & ssum_1_55; // @[Mul.scala 192:44]
  wire  _sum_T_685 = ssum_2_36 ^ cout_100; // @[Mul.scala 191:34]
  wire  ssum_0_104 = ssum_2_36 ^ cout_100 ^ scout_0_68; // @[Mul.scala 191:42]
  wire  scout_0_104 = ssum_2_36 & cout_100 | _sum_T_685 & scout_0_68; // @[Mul.scala 192:44]
  wire  ssum_1_77 = scout_1_54 ^ scout_2_35; // @[Mul.scala 206:34]
  wire  scout_1_77 = scout_1_54 & scout_2_35; // @[Mul.scala 207:34]
  wire  _sum_T_688 = sum_102 ^ ssum_0_70; // @[Mul.scala 191:34]
  wire  sum_180 = sum_102 ^ ssum_0_70 ^ ssum_1_56; // @[Mul.scala 191:42]
  wire  cout_180 = sum_102 & ssum_0_70 | _sum_T_688 & ssum_1_56; // @[Mul.scala 192:44]
  wire  _sum_T_690 = ssum_2_37 ^ cout_101; // @[Mul.scala 191:34]
  wire  ssum_0_105 = ssum_2_37 ^ cout_101 ^ scout_0_69; // @[Mul.scala 191:42]
  wire  scout_0_105 = ssum_2_37 & cout_101 | _sum_T_690 & scout_0_69; // @[Mul.scala 192:44]
  wire  ssum_1_78 = scout_1_55 ^ scout_2_36; // @[Mul.scala 206:34]
  wire  scout_1_78 = scout_1_55 & scout_2_36; // @[Mul.scala 207:34]
  wire  _sum_T_693 = sum_103 ^ ssum_0_71; // @[Mul.scala 191:34]
  wire  sum_181 = sum_103 ^ ssum_0_71 ^ ssum_1_57; // @[Mul.scala 191:42]
  wire  cout_181 = sum_103 & ssum_0_71 | _sum_T_693 & ssum_1_57; // @[Mul.scala 192:44]
  wire  _sum_T_695 = ssum_2_38 ^ cout_102; // @[Mul.scala 191:34]
  wire  ssum_0_106 = ssum_2_38 ^ cout_102 ^ scout_0_70; // @[Mul.scala 191:42]
  wire  scout_0_106 = ssum_2_38 & cout_102 | _sum_T_695 & scout_0_70; // @[Mul.scala 192:44]
  wire  ssum_1_79 = scout_1_56 ^ scout_2_37; // @[Mul.scala 206:34]
  wire  scout_1_79 = scout_1_56 & scout_2_37; // @[Mul.scala 207:34]
  wire  _sum_T_698 = sum_104 ^ ssum_0_72; // @[Mul.scala 191:34]
  wire  sum_182 = sum_104 ^ ssum_0_72 ^ ssum_1_58; // @[Mul.scala 191:42]
  wire  cout_182 = sum_104 & ssum_0_72 | _sum_T_698 & ssum_1_58; // @[Mul.scala 192:44]
  wire  _sum_T_700 = ssum_2_39 ^ cout_103; // @[Mul.scala 191:34]
  wire  ssum_0_107 = ssum_2_39 ^ cout_103 ^ scout_0_71; // @[Mul.scala 191:42]
  wire  scout_0_107 = ssum_2_39 & cout_103 | _sum_T_700 & scout_0_71; // @[Mul.scala 192:44]
  wire  ssum_1_80 = scout_1_57 ^ scout_2_38; // @[Mul.scala 206:34]
  wire  scout_1_80 = scout_1_57 & scout_2_38; // @[Mul.scala 207:34]
  wire  _sum_T_703 = sum_105 ^ ssum_0_73; // @[Mul.scala 191:34]
  wire  sum_183 = sum_105 ^ ssum_0_73 ^ ssum_1_59; // @[Mul.scala 191:42]
  wire  cout_183 = sum_105 & ssum_0_73 | _sum_T_703 & ssum_1_59; // @[Mul.scala 192:44]
  wire  _sum_T_705 = ssum_2_40 ^ cout_104; // @[Mul.scala 191:34]
  wire  ssum_0_108 = ssum_2_40 ^ cout_104 ^ scout_0_72; // @[Mul.scala 191:42]
  wire  scout_0_108 = ssum_2_40 & cout_104 | _sum_T_705 & scout_0_72; // @[Mul.scala 192:44]
  wire  ssum_1_81 = scout_1_58 ^ scout_2_39; // @[Mul.scala 206:34]
  wire  scout_1_81 = scout_1_58 & scout_2_39; // @[Mul.scala 207:34]
  wire  _sum_T_708 = sum_106 ^ ssum_0_74; // @[Mul.scala 191:34]
  wire  sum_184 = sum_106 ^ ssum_0_74 ^ ssum_1_60; // @[Mul.scala 191:42]
  wire  cout_184 = sum_106 & ssum_0_74 | _sum_T_708 & ssum_1_60; // @[Mul.scala 192:44]
  wire  _sum_T_710 = ssum_2_41 ^ cout_105; // @[Mul.scala 191:34]
  wire  ssum_0_109 = ssum_2_41 ^ cout_105 ^ scout_0_73; // @[Mul.scala 191:42]
  wire  scout_0_109 = ssum_2_41 & cout_105 | _sum_T_710 & scout_0_73; // @[Mul.scala 192:44]
  wire  ssum_1_82 = scout_1_59 ^ scout_2_40; // @[Mul.scala 206:34]
  wire  scout_1_82 = scout_1_59 & scout_2_40; // @[Mul.scala 207:34]
  wire  _sum_T_713 = sum_107 ^ ssum_0_75; // @[Mul.scala 191:34]
  wire  sum_185 = sum_107 ^ ssum_0_75 ^ ssum_1_61; // @[Mul.scala 191:42]
  wire  cout_185 = sum_107 & ssum_0_75 | _sum_T_713 & ssum_1_61; // @[Mul.scala 192:44]
  wire  _sum_T_715 = ssum_2_42 ^ cout_106; // @[Mul.scala 191:34]
  wire  ssum_0_110 = ssum_2_42 ^ cout_106 ^ scout_0_74; // @[Mul.scala 191:42]
  wire  scout_0_110 = ssum_2_42 & cout_106 | _sum_T_715 & scout_0_74; // @[Mul.scala 192:44]
  wire  ssum_1_83 = scout_1_60 ^ scout_2_41; // @[Mul.scala 206:34]
  wire  scout_1_83 = scout_1_60 & scout_2_41; // @[Mul.scala 207:34]
  wire  _sum_T_718 = sum_108 ^ ssum_0_76; // @[Mul.scala 191:34]
  wire  sum_186 = sum_108 ^ ssum_0_76 ^ ssum_1_62; // @[Mul.scala 191:42]
  wire  cout_186 = sum_108 & ssum_0_76 | _sum_T_718 & ssum_1_62; // @[Mul.scala 192:44]
  wire  ssum_0_111 = cout_107 ^ scout_0_75; // @[Mul.scala 206:34]
  wire  scout_0_111 = cout_107 & scout_0_75; // @[Mul.scala 207:34]
  wire  ssum_1_84 = scout_1_61 ^ scout_2_42; // @[Mul.scala 206:34]
  wire  scout_1_84 = scout_1_61 & scout_2_42; // @[Mul.scala 207:34]
  wire  _sum_T_722 = sum_109 ^ ssum_0_77; // @[Mul.scala 191:34]
  wire  sum_187 = sum_109 ^ ssum_0_77 ^ ssum_1_63; // @[Mul.scala 191:42]
  wire  cout_187 = sum_109 & ssum_0_77 | _sum_T_722 & ssum_1_63; // @[Mul.scala 192:44]
  wire  _sum_T_724 = cout_108 ^ scout_0_76; // @[Mul.scala 191:34]
  wire  ssum_0_112 = cout_108 ^ scout_0_76 ^ scout_1_62; // @[Mul.scala 191:42]
  wire  scout_0_112 = cout_108 & scout_0_76 | _sum_T_724 & scout_1_62; // @[Mul.scala 192:44]
  wire  _sum_T_726 = sum_110 ^ ssum_0_78; // @[Mul.scala 191:34]
  wire  sum_188 = sum_110 ^ ssum_0_78 ^ ssum_1_64; // @[Mul.scala 191:42]
  wire  cout_188 = sum_110 & ssum_0_78 | _sum_T_726 & ssum_1_64; // @[Mul.scala 192:44]
  wire  _sum_T_728 = cout_109 ^ scout_0_77; // @[Mul.scala 191:34]
  wire  ssum_0_113 = cout_109 ^ scout_0_77 ^ scout_1_63; // @[Mul.scala 191:42]
  wire  scout_0_113 = cout_109 & scout_0_77 | _sum_T_728 & scout_1_63; // @[Mul.scala 192:44]
  wire  _sum_T_730 = sum_111 ^ ssum_0_79; // @[Mul.scala 191:34]
  wire  sum_189 = sum_111 ^ ssum_0_79 ^ ssum_1_65; // @[Mul.scala 191:42]
  wire  cout_189 = sum_111 & ssum_0_79 | _sum_T_730 & ssum_1_65; // @[Mul.scala 192:44]
  wire  _sum_T_732 = cout_110 ^ scout_0_78; // @[Mul.scala 191:34]
  wire  ssum_0_114 = cout_110 ^ scout_0_78 ^ scout_1_64; // @[Mul.scala 191:42]
  wire  scout_0_114 = cout_110 & scout_0_78 | _sum_T_732 & scout_1_64; // @[Mul.scala 192:44]
  wire  _sum_T_734 = sum_112 ^ ssum_0_80; // @[Mul.scala 191:34]
  wire  sum_190 = sum_112 ^ ssum_0_80 ^ ssum_1_66; // @[Mul.scala 191:42]
  wire  cout_190 = sum_112 & ssum_0_80 | _sum_T_734 & ssum_1_66; // @[Mul.scala 192:44]
  wire  _sum_T_736 = cout_111 ^ scout_0_79; // @[Mul.scala 191:34]
  wire  ssum_0_115 = cout_111 ^ scout_0_79 ^ scout_1_65; // @[Mul.scala 191:42]
  wire  scout_0_115 = cout_111 & scout_0_79 | _sum_T_736 & scout_1_65; // @[Mul.scala 192:44]
  wire  _sum_T_738 = sum_113 ^ ssum_0_81; // @[Mul.scala 191:34]
  wire  sum_191 = sum_113 ^ ssum_0_81 ^ ssum_1_67; // @[Mul.scala 191:42]
  wire  cout_191 = sum_113 & ssum_0_81 | _sum_T_738 & ssum_1_67; // @[Mul.scala 192:44]
  wire  _sum_T_740 = cout_112 ^ scout_0_80; // @[Mul.scala 191:34]
  wire  ssum_0_116 = cout_112 ^ scout_0_80 ^ scout_1_66; // @[Mul.scala 191:42]
  wire  scout_0_116 = cout_112 & scout_0_80 | _sum_T_740 & scout_1_66; // @[Mul.scala 192:44]
  wire  _sum_T_742 = sum_114 ^ ssum_0_82; // @[Mul.scala 191:34]
  wire  sum_192 = sum_114 ^ ssum_0_82 ^ ssum_1_68; // @[Mul.scala 191:42]
  wire  cout_192 = sum_114 & ssum_0_82 | _sum_T_742 & ssum_1_68; // @[Mul.scala 192:44]
  wire  _sum_T_744 = cout_113 ^ scout_0_81; // @[Mul.scala 191:34]
  wire  ssum_0_117 = cout_113 ^ scout_0_81 ^ scout_1_67; // @[Mul.scala 191:42]
  wire  scout_0_117 = cout_113 & scout_0_81 | _sum_T_744 & scout_1_67; // @[Mul.scala 192:44]
  wire  _sum_T_746 = sum_115 ^ ssum_0_83; // @[Mul.scala 191:34]
  wire  sum_193 = sum_115 ^ ssum_0_83 ^ cout_114; // @[Mul.scala 191:42]
  wire  cout_193 = sum_115 & ssum_0_83 | _sum_T_746 & cout_114; // @[Mul.scala 192:44]
  wire  ssum_0_118 = scout_0_82 ^ scout_1_68; // @[Mul.scala 206:34]
  wire  scout_0_118 = scout_0_82 & scout_1_68; // @[Mul.scala 207:34]
  wire  sum_194 = sum_116 ^ ssum_0_84; // @[Mul.scala 206:34]
  wire  cout_194 = sum_116 & ssum_0_84; // @[Mul.scala 207:34]
  wire  sum_195 = cout_115 ^ scout_0_83; // @[Mul.scala 206:34]
  wire  cout_195 = cout_115 & scout_0_83; // @[Mul.scala 207:34]
  wire  sum_196 = sum_117 ^ ssum_0_85; // @[Mul.scala 206:34]
  wire  cout_196 = sum_117 & ssum_0_85; // @[Mul.scala 207:34]
  wire  sum_197 = cout_116 ^ scout_0_84; // @[Mul.scala 206:34]
  wire  cout_197 = cout_116 & scout_0_84; // @[Mul.scala 207:34]
  wire  sum_198 = sum_118 ^ ssum_0_86; // @[Mul.scala 206:34]
  wire  cout_198 = sum_118 & ssum_0_86; // @[Mul.scala 207:34]
  wire  sum_199 = cout_117 ^ scout_0_85; // @[Mul.scala 206:34]
  wire  cout_199 = cout_117 & scout_0_85; // @[Mul.scala 207:34]
  wire  sum_200 = sum_119 ^ ssum_0_87; // @[Mul.scala 206:34]
  wire  cout_200 = sum_119 & ssum_0_87; // @[Mul.scala 207:34]
  wire  sum_201 = cout_118 ^ scout_0_86; // @[Mul.scala 206:34]
  wire  cout_201 = cout_118 & scout_0_86; // @[Mul.scala 207:34]
  wire  sum_202 = sum_120 ^ ssum_0_88; // @[Mul.scala 206:34]
  wire  cout_202 = sum_120 & ssum_0_88; // @[Mul.scala 207:34]
  wire  sum_203 = cout_119 ^ scout_0_87; // @[Mul.scala 206:34]
  wire  cout_203 = cout_119 & scout_0_87; // @[Mul.scala 207:34]
  wire  sum_204 = sum_121 ^ sum_122; // @[Mul.scala 206:34]
  wire  cout_204 = sum_121 & sum_122; // @[Mul.scala 207:34]
  wire  sum_205 = cout_120 ^ scout_0_88; // @[Mul.scala 206:34]
  wire  cout_205 = cout_120 & scout_0_88; // @[Mul.scala 207:34]
  wire  sum_206 = sum_123 ^ sum_124; // @[Mul.scala 206:34]
  wire  cout_206 = sum_123 & sum_124; // @[Mul.scala 207:34]
  wire  sum_207 = cout_121 ^ cout_122; // @[Mul.scala 206:34]
  wire  cout_207 = cout_121 & cout_122; // @[Mul.scala 207:34]
  wire  sum_208 = sum_125 ^ sum_126; // @[Mul.scala 206:34]
  wire  cout_208 = sum_125 & sum_126; // @[Mul.scala 207:34]
  wire  sum_209 = cout_123 ^ cout_124; // @[Mul.scala 206:34]
  wire  cout_209 = cout_123 & cout_124; // @[Mul.scala 207:34]
  wire  sum_210 = sum_127 ^ sum_128; // @[Mul.scala 206:34]
  wire  cout_210 = sum_127 & sum_128; // @[Mul.scala 207:34]
  wire  sum_211 = cout_125 ^ cout_126; // @[Mul.scala 206:34]
  wire  cout_211 = cout_125 & cout_126; // @[Mul.scala 207:34]
  wire  sum_212 = sum_129 ^ sum_130; // @[Mul.scala 206:34]
  wire  cout_212 = sum_129 & sum_130; // @[Mul.scala 207:34]
  wire  sum_213 = cout_127 ^ cout_128; // @[Mul.scala 206:34]
  wire  cout_213 = cout_127 & cout_128; // @[Mul.scala 207:34]
  wire  _sum_T_769 = sum_131 ^ cout_129; // @[Mul.scala 191:34]
  wire  sum_214 = sum_131 ^ cout_129 ^ cout_130; // @[Mul.scala 191:42]
  wire  cout_214 = sum_131 & cout_129 | _sum_T_769 & cout_130; // @[Mul.scala 192:44]
  wire  sum_215 = sum_132 ^ cout_131; // @[Mul.scala 206:34]
  wire  cout_215 = sum_132 & cout_131; // @[Mul.scala 207:34]
  wire  sum_216 = sum_133 ^ cout_132; // @[Mul.scala 206:34]
  wire  cout_216 = sum_133 & cout_132; // @[Mul.scala 207:34]
  wire  sum_217 = sum_134 ^ cout_133; // @[Mul.scala 206:34]
  wire  cout_217 = sum_134 & cout_133; // @[Mul.scala 207:34]
  wire  sum_218 = sum_135 ^ cout_134; // @[Mul.scala 206:34]
  wire  cout_218 = sum_135 & cout_134; // @[Mul.scala 207:34]
  wire  sum_219 = tree_63_0 ^ cout_135; // @[Mul.scala 206:34]
  wire  sum_224 = sum_141 ^ cout_140; // @[Mul.scala 206:34]
  wire  cout_224 = sum_141 & cout_140; // @[Mul.scala 207:34]
  wire  sum_225 = sum_142 ^ cout_141; // @[Mul.scala 206:34]
  wire  cout_225 = sum_142 & cout_141; // @[Mul.scala 207:34]
  wire  sum_226 = sum_143 ^ cout_142; // @[Mul.scala 206:34]
  wire  cout_226 = sum_143 & cout_142; // @[Mul.scala 207:34]
  wire  _sum_T_783 = sum_144 ^ sum_145; // @[Mul.scala 191:34]
  wire  sum_227 = sum_144 ^ sum_145 ^ cout_143; // @[Mul.scala 191:42]
  wire  cout_227 = sum_144 & sum_145 | _sum_T_783 & cout_143; // @[Mul.scala 192:44]
  wire  sum_228 = sum_146 ^ sum_147; // @[Mul.scala 206:34]
  wire  cout_228 = sum_146 & sum_147; // @[Mul.scala 207:34]
  wire  sum_229 = cout_144 ^ cout_145; // @[Mul.scala 206:34]
  wire  cout_229 = cout_144 & cout_145; // @[Mul.scala 207:34]
  wire  sum_230 = sum_148 ^ sum_149; // @[Mul.scala 206:34]
  wire  cout_230 = sum_148 & sum_149; // @[Mul.scala 207:34]
  wire  sum_231 = cout_146 ^ cout_147; // @[Mul.scala 206:34]
  wire  cout_231 = cout_146 & cout_147; // @[Mul.scala 207:34]
  wire  sum_232 = sum_150 ^ sum_151; // @[Mul.scala 206:34]
  wire  cout_232 = sum_150 & sum_151; // @[Mul.scala 207:34]
  wire  sum_233 = cout_148 ^ cout_149; // @[Mul.scala 206:34]
  wire  cout_233 = cout_148 & cout_149; // @[Mul.scala 207:34]
  wire  sum_234 = sum_152 ^ sum_153; // @[Mul.scala 206:34]
  wire  cout_234 = sum_152 & sum_153; // @[Mul.scala 207:34]
  wire  sum_235 = cout_150 ^ cout_151; // @[Mul.scala 206:34]
  wire  cout_235 = cout_150 & cout_151; // @[Mul.scala 207:34]
  wire  sum_236 = sum_154 ^ sum_155; // @[Mul.scala 206:34]
  wire  cout_236 = sum_154 & sum_155; // @[Mul.scala 207:34]
  wire  sum_237 = cout_152 ^ cout_153; // @[Mul.scala 206:34]
  wire  cout_237 = cout_152 & cout_153; // @[Mul.scala 207:34]
  wire  sum_238 = sum_156 ^ sum_157; // @[Mul.scala 206:34]
  wire  cout_238 = sum_156 & sum_157; // @[Mul.scala 207:34]
  wire  sum_239 = cout_154 ^ cout_155; // @[Mul.scala 206:34]
  wire  cout_239 = cout_154 & cout_155; // @[Mul.scala 207:34]
  wire  sum_240 = sum_158 ^ sum_159; // @[Mul.scala 206:34]
  wire  cout_240 = sum_158 & sum_159; // @[Mul.scala 207:34]
  wire  sum_241 = cout_156 ^ cout_157; // @[Mul.scala 206:34]
  wire  cout_241 = cout_156 & cout_157; // @[Mul.scala 207:34]
  wire  sum_242 = sum_160 ^ sum_161; // @[Mul.scala 206:34]
  wire  cout_242 = sum_160 & sum_161; // @[Mul.scala 207:34]
  wire  sum_243 = cout_158 ^ cout_159; // @[Mul.scala 206:34]
  wire  cout_243 = cout_158 & cout_159; // @[Mul.scala 207:34]
  wire  sum_244 = sum_162 ^ sum_163; // @[Mul.scala 206:34]
  wire  cout_244 = sum_162 & sum_163; // @[Mul.scala 207:34]
  wire  sum_245 = cout_160 ^ cout_161; // @[Mul.scala 206:34]
  wire  cout_245 = cout_160 & cout_161; // @[Mul.scala 207:34]
  wire  sum_246 = sum_164 ^ ssum_0_89; // @[Mul.scala 206:34]
  wire  cout_246 = sum_164 & ssum_0_89; // @[Mul.scala 207:34]
  wire  sum_247 = cout_162 ^ cout_163; // @[Mul.scala 206:34]
  wire  cout_247 = cout_162 & cout_163; // @[Mul.scala 207:34]
  wire  sum_248 = sum_165 ^ ssum_0_90; // @[Mul.scala 206:34]
  wire  cout_248 = sum_165 & ssum_0_90; // @[Mul.scala 207:34]
  wire  sum_249 = cout_164 ^ scout_0_89; // @[Mul.scala 206:34]
  wire  cout_249 = cout_164 & scout_0_89; // @[Mul.scala 207:34]
  wire  sum_250 = sum_166 ^ ssum_0_91; // @[Mul.scala 206:34]
  wire  cout_250 = sum_166 & ssum_0_91; // @[Mul.scala 207:34]
  wire  sum_251 = cout_165 ^ scout_0_90; // @[Mul.scala 206:34]
  wire  cout_251 = cout_165 & scout_0_90; // @[Mul.scala 207:34]
  wire  sum_252 = sum_167 ^ ssum_0_92; // @[Mul.scala 206:34]
  wire  cout_252 = sum_167 & ssum_0_92; // @[Mul.scala 207:34]
  wire  sum_253 = cout_166 ^ scout_0_91; // @[Mul.scala 206:34]
  wire  cout_253 = cout_166 & scout_0_91; // @[Mul.scala 207:34]
  wire  sum_254 = sum_168 ^ ssum_0_93; // @[Mul.scala 206:34]
  wire  cout_254 = sum_168 & ssum_0_93; // @[Mul.scala 207:34]
  wire  sum_255 = cout_167 ^ scout_0_92; // @[Mul.scala 206:34]
  wire  cout_255 = cout_167 & scout_0_92; // @[Mul.scala 207:34]
  wire  sum_256 = sum_169 ^ ssum_0_94; // @[Mul.scala 206:34]
  wire  cout_256 = sum_169 & ssum_0_94; // @[Mul.scala 207:34]
  wire  sum_257 = cout_168 ^ scout_0_93; // @[Mul.scala 206:34]
  wire  cout_257 = cout_168 & scout_0_93; // @[Mul.scala 207:34]
  wire  sum_258 = sum_170 ^ ssum_0_95; // @[Mul.scala 206:34]
  wire  cout_258 = sum_170 & ssum_0_95; // @[Mul.scala 207:34]
  wire  sum_259 = cout_169 ^ scout_0_94; // @[Mul.scala 206:34]
  wire  cout_259 = cout_169 & scout_0_94; // @[Mul.scala 207:34]
  wire  _sum_T_817 = sum_171 ^ ssum_0_96; // @[Mul.scala 191:34]
  wire  sum_260 = sum_171 ^ ssum_0_96 ^ ssum_1_69; // @[Mul.scala 191:42]
  wire  cout_260 = sum_171 & ssum_0_96 | _sum_T_817 & ssum_1_69; // @[Mul.scala 192:44]
  wire  ssum_0_119 = cout_170 ^ scout_0_95; // @[Mul.scala 206:34]
  wire  scout_0_119 = cout_170 & scout_0_95; // @[Mul.scala 207:34]
  wire  _sum_T_820 = sum_172 ^ ssum_0_97; // @[Mul.scala 191:34]
  wire  sum_261 = sum_172 ^ ssum_0_97 ^ ssum_1_70; // @[Mul.scala 191:42]
  wire  cout_261 = sum_172 & ssum_0_97 | _sum_T_820 & ssum_1_70; // @[Mul.scala 192:44]
  wire  _sum_T_822 = cout_171 ^ scout_0_96; // @[Mul.scala 191:34]
  wire  ssum_0_120 = cout_171 ^ scout_0_96 ^ scout_1_69; // @[Mul.scala 191:42]
  wire  scout_0_120 = cout_171 & scout_0_96 | _sum_T_822 & scout_1_69; // @[Mul.scala 192:44]
  wire  _sum_T_824 = sum_173 ^ ssum_0_98; // @[Mul.scala 191:34]
  wire  sum_262 = sum_173 ^ ssum_0_98 ^ ssum_1_71; // @[Mul.scala 191:42]
  wire  cout_262 = sum_173 & ssum_0_98 | _sum_T_824 & ssum_1_71; // @[Mul.scala 192:44]
  wire  _sum_T_826 = cout_172 ^ scout_0_97; // @[Mul.scala 191:34]
  wire  ssum_0_121 = cout_172 ^ scout_0_97 ^ scout_1_70; // @[Mul.scala 191:42]
  wire  scout_0_121 = cout_172 & scout_0_97 | _sum_T_826 & scout_1_70; // @[Mul.scala 192:44]
  wire  _sum_T_828 = sum_174 ^ ssum_0_99; // @[Mul.scala 191:34]
  wire  sum_263 = sum_174 ^ ssum_0_99 ^ ssum_1_72; // @[Mul.scala 191:42]
  wire  cout_263 = sum_174 & ssum_0_99 | _sum_T_828 & ssum_1_72; // @[Mul.scala 192:44]
  wire  _sum_T_830 = cout_173 ^ scout_0_98; // @[Mul.scala 191:34]
  wire  ssum_0_122 = cout_173 ^ scout_0_98 ^ scout_1_71; // @[Mul.scala 191:42]
  wire  scout_0_122 = cout_173 & scout_0_98 | _sum_T_830 & scout_1_71; // @[Mul.scala 192:44]
  wire  _sum_T_832 = sum_175 ^ ssum_0_100; // @[Mul.scala 191:34]
  wire  sum_264 = sum_175 ^ ssum_0_100 ^ ssum_1_73; // @[Mul.scala 191:42]
  wire  cout_264 = sum_175 & ssum_0_100 | _sum_T_832 & ssum_1_73; // @[Mul.scala 192:44]
  wire  _sum_T_834 = cout_174 ^ scout_0_99; // @[Mul.scala 191:34]
  wire  ssum_0_123 = cout_174 ^ scout_0_99 ^ scout_1_72; // @[Mul.scala 191:42]
  wire  scout_0_123 = cout_174 & scout_0_99 | _sum_T_834 & scout_1_72; // @[Mul.scala 192:44]
  wire  _sum_T_836 = sum_176 ^ ssum_0_101; // @[Mul.scala 191:34]
  wire  sum_265 = sum_176 ^ ssum_0_101 ^ ssum_1_74; // @[Mul.scala 191:42]
  wire  cout_265 = sum_176 & ssum_0_101 | _sum_T_836 & ssum_1_74; // @[Mul.scala 192:44]
  wire  _sum_T_838 = cout_175 ^ scout_0_100; // @[Mul.scala 191:34]
  wire  ssum_0_124 = cout_175 ^ scout_0_100 ^ scout_1_73; // @[Mul.scala 191:42]
  wire  scout_0_124 = cout_175 & scout_0_100 | _sum_T_838 & scout_1_73; // @[Mul.scala 192:44]
  wire  _sum_T_840 = sum_177 ^ ssum_0_102; // @[Mul.scala 191:34]
  wire  sum_266 = sum_177 ^ ssum_0_102 ^ ssum_1_75; // @[Mul.scala 191:42]
  wire  cout_266 = sum_177 & ssum_0_102 | _sum_T_840 & ssum_1_75; // @[Mul.scala 192:44]
  wire  _sum_T_842 = cout_176 ^ scout_0_101; // @[Mul.scala 191:34]
  wire  ssum_0_125 = cout_176 ^ scout_0_101 ^ scout_1_74; // @[Mul.scala 191:42]
  wire  scout_0_125 = cout_176 & scout_0_101 | _sum_T_842 & scout_1_74; // @[Mul.scala 192:44]
  wire  _sum_T_844 = sum_178 ^ ssum_0_103; // @[Mul.scala 191:34]
  wire  sum_267 = sum_178 ^ ssum_0_103 ^ ssum_1_76; // @[Mul.scala 191:42]
  wire  cout_267 = sum_178 & ssum_0_103 | _sum_T_844 & ssum_1_76; // @[Mul.scala 192:44]
  wire  _sum_T_846 = cout_177 ^ scout_0_102; // @[Mul.scala 191:34]
  wire  ssum_0_126 = cout_177 ^ scout_0_102 ^ scout_1_75; // @[Mul.scala 191:42]
  wire  scout_0_126 = cout_177 & scout_0_102 | _sum_T_846 & scout_1_75; // @[Mul.scala 192:44]
  wire  _sum_T_848 = sum_179 ^ ssum_0_104; // @[Mul.scala 191:34]
  wire  sum_268 = sum_179 ^ ssum_0_104 ^ ssum_1_77; // @[Mul.scala 191:42]
  wire  cout_268 = sum_179 & ssum_0_104 | _sum_T_848 & ssum_1_77; // @[Mul.scala 192:44]
  wire  _sum_T_850 = cout_178 ^ scout_0_103; // @[Mul.scala 191:34]
  wire  ssum_0_127 = cout_178 ^ scout_0_103 ^ scout_1_76; // @[Mul.scala 191:42]
  wire  scout_0_127 = cout_178 & scout_0_103 | _sum_T_850 & scout_1_76; // @[Mul.scala 192:44]
  wire  _sum_T_852 = sum_180 ^ ssum_0_105; // @[Mul.scala 191:34]
  wire  sum_269 = sum_180 ^ ssum_0_105 ^ ssum_1_78; // @[Mul.scala 191:42]
  wire  cout_269 = sum_180 & ssum_0_105 | _sum_T_852 & ssum_1_78; // @[Mul.scala 192:44]
  wire  _sum_T_854 = cout_179 ^ scout_0_104; // @[Mul.scala 191:34]
  wire  ssum_0_128 = cout_179 ^ scout_0_104 ^ scout_1_77; // @[Mul.scala 191:42]
  wire  scout_0_128 = cout_179 & scout_0_104 | _sum_T_854 & scout_1_77; // @[Mul.scala 192:44]
  wire  _sum_T_856 = sum_181 ^ ssum_0_106; // @[Mul.scala 191:34]
  wire  sum_270 = sum_181 ^ ssum_0_106 ^ ssum_1_79; // @[Mul.scala 191:42]
  wire  cout_270 = sum_181 & ssum_0_106 | _sum_T_856 & ssum_1_79; // @[Mul.scala 192:44]
  wire  _sum_T_858 = cout_180 ^ scout_0_105; // @[Mul.scala 191:34]
  wire  ssum_0_129 = cout_180 ^ scout_0_105 ^ scout_1_78; // @[Mul.scala 191:42]
  wire  scout_0_129 = cout_180 & scout_0_105 | _sum_T_858 & scout_1_78; // @[Mul.scala 192:44]
  wire  _sum_T_860 = sum_182 ^ ssum_0_107; // @[Mul.scala 191:34]
  wire  sum_271 = sum_182 ^ ssum_0_107 ^ ssum_1_80; // @[Mul.scala 191:42]
  wire  cout_271 = sum_182 & ssum_0_107 | _sum_T_860 & ssum_1_80; // @[Mul.scala 192:44]
  wire  _sum_T_862 = cout_181 ^ scout_0_106; // @[Mul.scala 191:34]
  wire  ssum_0_130 = cout_181 ^ scout_0_106 ^ scout_1_79; // @[Mul.scala 191:42]
  wire  scout_0_130 = cout_181 & scout_0_106 | _sum_T_862 & scout_1_79; // @[Mul.scala 192:44]
  wire  _sum_T_864 = sum_183 ^ ssum_0_108; // @[Mul.scala 191:34]
  wire  sum_272 = sum_183 ^ ssum_0_108 ^ ssum_1_81; // @[Mul.scala 191:42]
  wire  cout_272 = sum_183 & ssum_0_108 | _sum_T_864 & ssum_1_81; // @[Mul.scala 192:44]
  wire  _sum_T_866 = cout_182 ^ scout_0_107; // @[Mul.scala 191:34]
  wire  ssum_0_131 = cout_182 ^ scout_0_107 ^ scout_1_80; // @[Mul.scala 191:42]
  wire  scout_0_131 = cout_182 & scout_0_107 | _sum_T_866 & scout_1_80; // @[Mul.scala 192:44]
  wire  _sum_T_868 = sum_184 ^ ssum_0_109; // @[Mul.scala 191:34]
  wire  sum_273 = sum_184 ^ ssum_0_109 ^ ssum_1_82; // @[Mul.scala 191:42]
  wire  cout_273 = sum_184 & ssum_0_109 | _sum_T_868 & ssum_1_82; // @[Mul.scala 192:44]
  wire  _sum_T_870 = cout_183 ^ scout_0_108; // @[Mul.scala 191:34]
  wire  ssum_0_132 = cout_183 ^ scout_0_108 ^ scout_1_81; // @[Mul.scala 191:42]
  wire  scout_0_132 = cout_183 & scout_0_108 | _sum_T_870 & scout_1_81; // @[Mul.scala 192:44]
  wire  _sum_T_872 = sum_185 ^ ssum_0_110; // @[Mul.scala 191:34]
  wire  sum_274 = sum_185 ^ ssum_0_110 ^ ssum_1_83; // @[Mul.scala 191:42]
  wire  cout_274 = sum_185 & ssum_0_110 | _sum_T_872 & ssum_1_83; // @[Mul.scala 192:44]
  wire  _sum_T_874 = cout_184 ^ scout_0_109; // @[Mul.scala 191:34]
  wire  ssum_0_133 = cout_184 ^ scout_0_109 ^ scout_1_82; // @[Mul.scala 191:42]
  wire  scout_0_133 = cout_184 & scout_0_109 | _sum_T_874 & scout_1_82; // @[Mul.scala 192:44]
  wire  _sum_T_876 = sum_186 ^ ssum_0_111; // @[Mul.scala 191:34]
  wire  sum_275 = sum_186 ^ ssum_0_111 ^ ssum_1_84; // @[Mul.scala 191:42]
  wire  cout_275 = sum_186 & ssum_0_111 | _sum_T_876 & ssum_1_84; // @[Mul.scala 192:44]
  wire  _sum_T_878 = cout_185 ^ scout_0_110; // @[Mul.scala 191:34]
  wire  ssum_0_134 = cout_185 ^ scout_0_110 ^ scout_1_83; // @[Mul.scala 191:42]
  wire  scout_0_134 = cout_185 & scout_0_110 | _sum_T_878 & scout_1_83; // @[Mul.scala 192:44]
  wire  _sum_T_880 = sum_187 ^ ssum_0_112; // @[Mul.scala 191:34]
  wire  sum_276 = sum_187 ^ ssum_0_112 ^ cout_186; // @[Mul.scala 191:42]
  wire  cout_276 = sum_187 & ssum_0_112 | _sum_T_880 & cout_186; // @[Mul.scala 192:44]
  wire  ssum_0_135 = scout_0_111 ^ scout_1_84; // @[Mul.scala 206:34]
  wire  scout_0_135 = scout_0_111 & scout_1_84; // @[Mul.scala 207:34]
  wire  sum_277 = sum_188 ^ ssum_0_113; // @[Mul.scala 206:34]
  wire  cout_277 = sum_188 & ssum_0_113; // @[Mul.scala 207:34]
  wire  sum_278 = cout_187 ^ scout_0_112; // @[Mul.scala 206:34]
  wire  cout_278 = cout_187 & scout_0_112; // @[Mul.scala 207:34]
  wire  sum_279 = sum_189 ^ ssum_0_114; // @[Mul.scala 206:34]
  wire  cout_279 = sum_189 & ssum_0_114; // @[Mul.scala 207:34]
  wire  sum_280 = cout_188 ^ scout_0_113; // @[Mul.scala 206:34]
  wire  cout_280 = cout_188 & scout_0_113; // @[Mul.scala 207:34]
  wire  sum_281 = sum_190 ^ ssum_0_115; // @[Mul.scala 206:34]
  wire  cout_281 = sum_190 & ssum_0_115; // @[Mul.scala 207:34]
  wire  sum_282 = cout_189 ^ scout_0_114; // @[Mul.scala 206:34]
  wire  cout_282 = cout_189 & scout_0_114; // @[Mul.scala 207:34]
  wire  sum_283 = sum_191 ^ ssum_0_116; // @[Mul.scala 206:34]
  wire  cout_283 = sum_191 & ssum_0_116; // @[Mul.scala 207:34]
  wire  sum_284 = cout_190 ^ scout_0_115; // @[Mul.scala 206:34]
  wire  cout_284 = cout_190 & scout_0_115; // @[Mul.scala 207:34]
  wire  sum_285 = sum_192 ^ ssum_0_117; // @[Mul.scala 206:34]
  wire  cout_285 = sum_192 & ssum_0_117; // @[Mul.scala 207:34]
  wire  sum_286 = cout_191 ^ scout_0_116; // @[Mul.scala 206:34]
  wire  cout_286 = cout_191 & scout_0_116; // @[Mul.scala 207:34]
  wire  sum_287 = sum_193 ^ ssum_0_118; // @[Mul.scala 206:34]
  wire  cout_287 = sum_193 & ssum_0_118; // @[Mul.scala 207:34]
  wire  sum_288 = cout_192 ^ scout_0_117; // @[Mul.scala 206:34]
  wire  cout_288 = cout_192 & scout_0_117; // @[Mul.scala 207:34]
  wire  sum_289 = sum_194 ^ sum_195; // @[Mul.scala 206:34]
  wire  cout_289 = sum_194 & sum_195; // @[Mul.scala 207:34]
  wire  sum_290 = cout_193 ^ scout_0_118; // @[Mul.scala 206:34]
  wire  cout_290 = cout_193 & scout_0_118; // @[Mul.scala 207:34]
  wire  sum_291 = sum_196 ^ sum_197; // @[Mul.scala 206:34]
  wire  cout_291 = sum_196 & sum_197; // @[Mul.scala 207:34]
  wire  sum_292 = cout_194 ^ cout_195; // @[Mul.scala 206:34]
  wire  cout_292 = cout_194 & cout_195; // @[Mul.scala 207:34]
  wire  sum_293 = sum_198 ^ sum_199; // @[Mul.scala 206:34]
  wire  cout_293 = sum_198 & sum_199; // @[Mul.scala 207:34]
  wire  sum_294 = cout_196 ^ cout_197; // @[Mul.scala 206:34]
  wire  cout_294 = cout_196 & cout_197; // @[Mul.scala 207:34]
  wire  sum_295 = sum_200 ^ sum_201; // @[Mul.scala 206:34]
  wire  cout_295 = sum_200 & sum_201; // @[Mul.scala 207:34]
  wire  sum_296 = cout_198 ^ cout_199; // @[Mul.scala 206:34]
  wire  cout_296 = cout_198 & cout_199; // @[Mul.scala 207:34]
  wire  sum_297 = sum_202 ^ sum_203; // @[Mul.scala 206:34]
  wire  cout_297 = sum_202 & sum_203; // @[Mul.scala 207:34]
  wire  sum_298 = cout_200 ^ cout_201; // @[Mul.scala 206:34]
  wire  cout_298 = cout_200 & cout_201; // @[Mul.scala 207:34]
  wire  sum_299 = sum_204 ^ sum_205; // @[Mul.scala 206:34]
  wire  cout_299 = sum_204 & sum_205; // @[Mul.scala 207:34]
  wire  sum_300 = cout_202 ^ cout_203; // @[Mul.scala 206:34]
  wire  cout_300 = cout_202 & cout_203; // @[Mul.scala 207:34]
  wire  sum_301 = sum_206 ^ sum_207; // @[Mul.scala 206:34]
  wire  cout_301 = sum_206 & sum_207; // @[Mul.scala 207:34]
  wire  sum_302 = cout_204 ^ cout_205; // @[Mul.scala 206:34]
  wire  cout_302 = cout_204 & cout_205; // @[Mul.scala 207:34]
  wire  sum_303 = sum_208 ^ sum_209; // @[Mul.scala 206:34]
  wire  cout_303 = sum_208 & sum_209; // @[Mul.scala 207:34]
  wire  sum_304 = cout_206 ^ cout_207; // @[Mul.scala 206:34]
  wire  cout_304 = cout_206 & cout_207; // @[Mul.scala 207:34]
  wire  sum_305 = sum_210 ^ sum_211; // @[Mul.scala 206:34]
  wire  cout_305 = sum_210 & sum_211; // @[Mul.scala 207:34]
  wire  sum_306 = cout_208 ^ cout_209; // @[Mul.scala 206:34]
  wire  cout_306 = cout_208 & cout_209; // @[Mul.scala 207:34]
  wire  sum_307 = sum_212 ^ sum_213; // @[Mul.scala 206:34]
  wire  cout_307 = sum_212 & sum_213; // @[Mul.scala 207:34]
  wire  sum_308 = cout_210 ^ cout_211; // @[Mul.scala 206:34]
  wire  cout_308 = cout_210 & cout_211; // @[Mul.scala 207:34]
  wire  _sum_T_915 = sum_214 ^ cout_212; // @[Mul.scala 191:34]
  wire  sum_309 = sum_214 ^ cout_212 ^ cout_213; // @[Mul.scala 191:42]
  wire  cout_309 = sum_214 & cout_212 | _sum_T_915 & cout_213; // @[Mul.scala 192:44]
  wire  sum_310 = sum_215 ^ cout_214; // @[Mul.scala 206:34]
  wire  cout_310 = sum_215 & cout_214; // @[Mul.scala 207:34]
  wire  sum_311 = sum_216 ^ cout_215; // @[Mul.scala 206:34]
  wire  cout_311 = sum_216 & cout_215; // @[Mul.scala 207:34]
  wire  sum_312 = sum_217 ^ cout_216; // @[Mul.scala 206:34]
  wire  cout_312 = sum_217 & cout_216; // @[Mul.scala 207:34]
  wire  sum_313 = sum_218 ^ cout_217; // @[Mul.scala 206:34]
  wire  cout_313 = sum_218 & cout_217; // @[Mul.scala 207:34]
  wire  sum_314 = sum_219 ^ cout_218; // @[Mul.scala 206:34]
  wire  sum_320 = sum_225 ^ cout_224; // @[Mul.scala 206:34]
  wire  cout_320 = sum_225 & cout_224; // @[Mul.scala 207:34]
  wire  sum_321 = sum_226 ^ cout_225; // @[Mul.scala 206:34]
  wire  cout_321 = sum_226 & cout_225; // @[Mul.scala 207:34]
  wire  sum_322 = sum_227 ^ cout_226; // @[Mul.scala 206:34]
  wire  cout_322 = sum_227 & cout_226; // @[Mul.scala 207:34]
  wire  _sum_T_930 = sum_228 ^ sum_229; // @[Mul.scala 191:34]
  wire  sum_323 = sum_228 ^ sum_229 ^ cout_227; // @[Mul.scala 191:42]
  wire  cout_323 = sum_228 & sum_229 | _sum_T_930 & cout_227; // @[Mul.scala 192:44]
  wire  sum_324 = sum_230 ^ sum_231; // @[Mul.scala 206:34]
  wire  cout_324 = sum_230 & sum_231; // @[Mul.scala 207:34]
  wire  sum_325 = cout_228 ^ cout_229; // @[Mul.scala 206:34]
  wire  cout_325 = cout_228 & cout_229; // @[Mul.scala 207:34]
  wire  sum_326 = sum_232 ^ sum_233; // @[Mul.scala 206:34]
  wire  cout_326 = sum_232 & sum_233; // @[Mul.scala 207:34]
  wire  sum_327 = cout_230 ^ cout_231; // @[Mul.scala 206:34]
  wire  cout_327 = cout_230 & cout_231; // @[Mul.scala 207:34]
  wire  sum_328 = sum_234 ^ sum_235; // @[Mul.scala 206:34]
  wire  cout_328 = sum_234 & sum_235; // @[Mul.scala 207:34]
  wire  sum_329 = cout_232 ^ cout_233; // @[Mul.scala 206:34]
  wire  cout_329 = cout_232 & cout_233; // @[Mul.scala 207:34]
  wire  sum_330 = sum_236 ^ sum_237; // @[Mul.scala 206:34]
  wire  cout_330 = sum_236 & sum_237; // @[Mul.scala 207:34]
  wire  sum_331 = cout_234 ^ cout_235; // @[Mul.scala 206:34]
  wire  cout_331 = cout_234 & cout_235; // @[Mul.scala 207:34]
  wire  sum_332 = sum_238 ^ sum_239; // @[Mul.scala 206:34]
  wire  cout_332 = sum_238 & sum_239; // @[Mul.scala 207:34]
  wire  sum_333 = cout_236 ^ cout_237; // @[Mul.scala 206:34]
  wire  cout_333 = cout_236 & cout_237; // @[Mul.scala 207:34]
  wire  sum_334 = sum_240 ^ sum_241; // @[Mul.scala 206:34]
  wire  cout_334 = sum_240 & sum_241; // @[Mul.scala 207:34]
  wire  sum_335 = cout_238 ^ cout_239; // @[Mul.scala 206:34]
  wire  cout_335 = cout_238 & cout_239; // @[Mul.scala 207:34]
  wire  sum_336 = sum_242 ^ sum_243; // @[Mul.scala 206:34]
  wire  cout_336 = sum_242 & sum_243; // @[Mul.scala 207:34]
  wire  sum_337 = cout_240 ^ cout_241; // @[Mul.scala 206:34]
  wire  cout_337 = cout_240 & cout_241; // @[Mul.scala 207:34]
  wire  sum_338 = sum_244 ^ sum_245; // @[Mul.scala 206:34]
  wire  cout_338 = sum_244 & sum_245; // @[Mul.scala 207:34]
  wire  sum_339 = cout_242 ^ cout_243; // @[Mul.scala 206:34]
  wire  cout_339 = cout_242 & cout_243; // @[Mul.scala 207:34]
  wire  sum_340 = sum_246 ^ sum_247; // @[Mul.scala 206:34]
  wire  cout_340 = sum_246 & sum_247; // @[Mul.scala 207:34]
  wire  sum_341 = cout_244 ^ cout_245; // @[Mul.scala 206:34]
  wire  cout_341 = cout_244 & cout_245; // @[Mul.scala 207:34]
  wire  sum_342 = sum_248 ^ sum_249; // @[Mul.scala 206:34]
  wire  cout_342 = sum_248 & sum_249; // @[Mul.scala 207:34]
  wire  sum_343 = cout_246 ^ cout_247; // @[Mul.scala 206:34]
  wire  cout_343 = cout_246 & cout_247; // @[Mul.scala 207:34]
  wire  sum_344 = sum_250 ^ sum_251; // @[Mul.scala 206:34]
  wire  cout_344 = sum_250 & sum_251; // @[Mul.scala 207:34]
  wire  sum_345 = cout_248 ^ cout_249; // @[Mul.scala 206:34]
  wire  cout_345 = cout_248 & cout_249; // @[Mul.scala 207:34]
  wire  sum_346 = sum_252 ^ sum_253; // @[Mul.scala 206:34]
  wire  cout_346 = sum_252 & sum_253; // @[Mul.scala 207:34]
  wire  sum_347 = cout_250 ^ cout_251; // @[Mul.scala 206:34]
  wire  cout_347 = cout_250 & cout_251; // @[Mul.scala 207:34]
  wire  sum_348 = sum_254 ^ sum_255; // @[Mul.scala 206:34]
  wire  cout_348 = sum_254 & sum_255; // @[Mul.scala 207:34]
  wire  sum_349 = cout_252 ^ cout_253; // @[Mul.scala 206:34]
  wire  cout_349 = cout_252 & cout_253; // @[Mul.scala 207:34]
  wire  sum_350 = sum_256 ^ sum_257; // @[Mul.scala 206:34]
  wire  cout_350 = sum_256 & sum_257; // @[Mul.scala 207:34]
  wire  sum_351 = cout_254 ^ cout_255; // @[Mul.scala 206:34]
  wire  cout_351 = cout_254 & cout_255; // @[Mul.scala 207:34]
  wire  sum_352 = sum_258 ^ sum_259; // @[Mul.scala 206:34]
  wire  cout_352 = sum_258 & sum_259; // @[Mul.scala 207:34]
  wire  sum_353 = cout_256 ^ cout_257; // @[Mul.scala 206:34]
  wire  cout_353 = cout_256 & cout_257; // @[Mul.scala 207:34]
  wire  sum_354 = sum_260 ^ ssum_0_119; // @[Mul.scala 206:34]
  wire  cout_354 = sum_260 & ssum_0_119; // @[Mul.scala 207:34]
  wire  sum_355 = cout_258 ^ cout_259; // @[Mul.scala 206:34]
  wire  cout_355 = cout_258 & cout_259; // @[Mul.scala 207:34]
  wire  sum_356 = sum_261 ^ ssum_0_120; // @[Mul.scala 206:34]
  wire  cout_356 = sum_261 & ssum_0_120; // @[Mul.scala 207:34]
  wire  sum_357 = cout_260 ^ scout_0_119; // @[Mul.scala 206:34]
  wire  cout_357 = cout_260 & scout_0_119; // @[Mul.scala 207:34]
  wire  sum_358 = sum_262 ^ ssum_0_121; // @[Mul.scala 206:34]
  wire  cout_358 = sum_262 & ssum_0_121; // @[Mul.scala 207:34]
  wire  sum_359 = cout_261 ^ scout_0_120; // @[Mul.scala 206:34]
  wire  cout_359 = cout_261 & scout_0_120; // @[Mul.scala 207:34]
  wire  sum_360 = sum_263 ^ ssum_0_122; // @[Mul.scala 206:34]
  wire  cout_360 = sum_263 & ssum_0_122; // @[Mul.scala 207:34]
  wire  sum_361 = cout_262 ^ scout_0_121; // @[Mul.scala 206:34]
  wire  cout_361 = cout_262 & scout_0_121; // @[Mul.scala 207:34]
  wire  sum_362 = sum_264 ^ ssum_0_123; // @[Mul.scala 206:34]
  wire  cout_362 = sum_264 & ssum_0_123; // @[Mul.scala 207:34]
  wire  sum_363 = cout_263 ^ scout_0_122; // @[Mul.scala 206:34]
  wire  cout_363 = cout_263 & scout_0_122; // @[Mul.scala 207:34]
  wire  sum_364 = sum_265 ^ ssum_0_124; // @[Mul.scala 206:34]
  wire  cout_364 = sum_265 & ssum_0_124; // @[Mul.scala 207:34]
  wire  sum_365 = cout_264 ^ scout_0_123; // @[Mul.scala 206:34]
  wire  cout_365 = cout_264 & scout_0_123; // @[Mul.scala 207:34]
  wire  sum_366 = sum_266 ^ ssum_0_125; // @[Mul.scala 206:34]
  wire  cout_366 = sum_266 & ssum_0_125; // @[Mul.scala 207:34]
  wire  sum_367 = cout_265 ^ scout_0_124; // @[Mul.scala 206:34]
  wire  cout_367 = cout_265 & scout_0_124; // @[Mul.scala 207:34]
  wire  sum_368 = sum_267 ^ ssum_0_126; // @[Mul.scala 206:34]
  wire  cout_368 = sum_267 & ssum_0_126; // @[Mul.scala 207:34]
  wire  sum_369 = cout_266 ^ scout_0_125; // @[Mul.scala 206:34]
  wire  cout_369 = cout_266 & scout_0_125; // @[Mul.scala 207:34]
  wire  sum_370 = sum_268 ^ ssum_0_127; // @[Mul.scala 206:34]
  wire  cout_370 = sum_268 & ssum_0_127; // @[Mul.scala 207:34]
  wire  sum_371 = cout_267 ^ scout_0_126; // @[Mul.scala 206:34]
  wire  cout_371 = cout_267 & scout_0_126; // @[Mul.scala 207:34]
  wire  sum_372 = sum_269 ^ ssum_0_128; // @[Mul.scala 206:34]
  wire  cout_372 = sum_269 & ssum_0_128; // @[Mul.scala 207:34]
  wire  sum_373 = cout_268 ^ scout_0_127; // @[Mul.scala 206:34]
  wire  cout_373 = cout_268 & scout_0_127; // @[Mul.scala 207:34]
  wire  sum_374 = sum_270 ^ ssum_0_129; // @[Mul.scala 206:34]
  wire  cout_374 = sum_270 & ssum_0_129; // @[Mul.scala 207:34]
  wire  sum_375 = cout_269 ^ scout_0_128; // @[Mul.scala 206:34]
  wire  cout_375 = cout_269 & scout_0_128; // @[Mul.scala 207:34]
  wire  sum_376 = sum_271 ^ ssum_0_130; // @[Mul.scala 206:34]
  wire  cout_376 = sum_271 & ssum_0_130; // @[Mul.scala 207:34]
  wire  sum_377 = cout_270 ^ scout_0_129; // @[Mul.scala 206:34]
  wire  cout_377 = cout_270 & scout_0_129; // @[Mul.scala 207:34]
  wire  sum_378 = sum_272 ^ ssum_0_131; // @[Mul.scala 206:34]
  wire  cout_378 = sum_272 & ssum_0_131; // @[Mul.scala 207:34]
  wire  sum_379 = cout_271 ^ scout_0_130; // @[Mul.scala 206:34]
  wire  cout_379 = cout_271 & scout_0_130; // @[Mul.scala 207:34]
  wire  sum_380 = sum_273 ^ ssum_0_132; // @[Mul.scala 206:34]
  wire  cout_380 = sum_273 & ssum_0_132; // @[Mul.scala 207:34]
  wire  sum_381 = cout_272 ^ scout_0_131; // @[Mul.scala 206:34]
  wire  cout_381 = cout_272 & scout_0_131; // @[Mul.scala 207:34]
  wire  sum_382 = sum_274 ^ ssum_0_133; // @[Mul.scala 206:34]
  wire  cout_382 = sum_274 & ssum_0_133; // @[Mul.scala 207:34]
  wire  sum_383 = cout_273 ^ scout_0_132; // @[Mul.scala 206:34]
  wire  cout_383 = cout_273 & scout_0_132; // @[Mul.scala 207:34]
  wire  sum_384 = sum_275 ^ ssum_0_134; // @[Mul.scala 206:34]
  wire  cout_384 = sum_275 & ssum_0_134; // @[Mul.scala 207:34]
  wire  sum_385 = cout_274 ^ scout_0_133; // @[Mul.scala 206:34]
  wire  cout_385 = cout_274 & scout_0_133; // @[Mul.scala 207:34]
  wire  sum_386 = sum_276 ^ ssum_0_135; // @[Mul.scala 206:34]
  wire  cout_386 = sum_276 & ssum_0_135; // @[Mul.scala 207:34]
  wire  sum_387 = cout_275 ^ scout_0_134; // @[Mul.scala 206:34]
  wire  cout_387 = cout_275 & scout_0_134; // @[Mul.scala 207:34]
  wire  sum_388 = sum_277 ^ sum_278; // @[Mul.scala 206:34]
  wire  cout_388 = sum_277 & sum_278; // @[Mul.scala 207:34]
  wire  sum_389 = cout_276 ^ scout_0_135; // @[Mul.scala 206:34]
  wire  cout_389 = cout_276 & scout_0_135; // @[Mul.scala 207:34]
  wire  sum_390 = sum_279 ^ sum_280; // @[Mul.scala 206:34]
  wire  cout_390 = sum_279 & sum_280; // @[Mul.scala 207:34]
  wire  sum_391 = cout_277 ^ cout_278; // @[Mul.scala 206:34]
  wire  cout_391 = cout_277 & cout_278; // @[Mul.scala 207:34]
  wire  sum_392 = sum_281 ^ sum_282; // @[Mul.scala 206:34]
  wire  cout_392 = sum_281 & sum_282; // @[Mul.scala 207:34]
  wire  sum_393 = cout_279 ^ cout_280; // @[Mul.scala 206:34]
  wire  cout_393 = cout_279 & cout_280; // @[Mul.scala 207:34]
  wire  sum_394 = sum_283 ^ sum_284; // @[Mul.scala 206:34]
  wire  cout_394 = sum_283 & sum_284; // @[Mul.scala 207:34]
  wire  sum_395 = cout_281 ^ cout_282; // @[Mul.scala 206:34]
  wire  cout_395 = cout_281 & cout_282; // @[Mul.scala 207:34]
  wire  sum_396 = sum_285 ^ sum_286; // @[Mul.scala 206:34]
  wire  cout_396 = sum_285 & sum_286; // @[Mul.scala 207:34]
  wire  sum_397 = cout_283 ^ cout_284; // @[Mul.scala 206:34]
  wire  cout_397 = cout_283 & cout_284; // @[Mul.scala 207:34]
  wire  sum_398 = sum_287 ^ sum_288; // @[Mul.scala 206:34]
  wire  cout_398 = sum_287 & sum_288; // @[Mul.scala 207:34]
  wire  sum_399 = cout_285 ^ cout_286; // @[Mul.scala 206:34]
  wire  cout_399 = cout_285 & cout_286; // @[Mul.scala 207:34]
  wire  sum_400 = sum_289 ^ sum_290; // @[Mul.scala 206:34]
  wire  cout_400 = sum_289 & sum_290; // @[Mul.scala 207:34]
  wire  sum_401 = cout_287 ^ cout_288; // @[Mul.scala 206:34]
  wire  cout_401 = cout_287 & cout_288; // @[Mul.scala 207:34]
  wire  sum_402 = sum_291 ^ sum_292; // @[Mul.scala 206:34]
  wire  cout_402 = sum_291 & sum_292; // @[Mul.scala 207:34]
  wire  sum_403 = cout_289 ^ cout_290; // @[Mul.scala 206:34]
  wire  cout_403 = cout_289 & cout_290; // @[Mul.scala 207:34]
  wire  sum_404 = sum_293 ^ sum_294; // @[Mul.scala 206:34]
  wire  cout_404 = sum_293 & sum_294; // @[Mul.scala 207:34]
  wire  sum_405 = cout_291 ^ cout_292; // @[Mul.scala 206:34]
  wire  cout_405 = cout_291 & cout_292; // @[Mul.scala 207:34]
  wire  sum_406 = sum_295 ^ sum_296; // @[Mul.scala 206:34]
  wire  cout_406 = sum_295 & sum_296; // @[Mul.scala 207:34]
  wire  sum_407 = cout_293 ^ cout_294; // @[Mul.scala 206:34]
  wire  cout_407 = cout_293 & cout_294; // @[Mul.scala 207:34]
  wire  sum_408 = sum_297 ^ sum_298; // @[Mul.scala 206:34]
  wire  cout_408 = sum_297 & sum_298; // @[Mul.scala 207:34]
  wire  sum_409 = cout_295 ^ cout_296; // @[Mul.scala 206:34]
  wire  cout_409 = cout_295 & cout_296; // @[Mul.scala 207:34]
  wire  sum_410 = sum_299 ^ sum_300; // @[Mul.scala 206:34]
  wire  cout_410 = sum_299 & sum_300; // @[Mul.scala 207:34]
  wire  sum_411 = cout_297 ^ cout_298; // @[Mul.scala 206:34]
  wire  cout_411 = cout_297 & cout_298; // @[Mul.scala 207:34]
  wire  sum_412 = sum_301 ^ sum_302; // @[Mul.scala 206:34]
  wire  cout_412 = sum_301 & sum_302; // @[Mul.scala 207:34]
  wire  sum_413 = cout_299 ^ cout_300; // @[Mul.scala 206:34]
  wire  cout_413 = cout_299 & cout_300; // @[Mul.scala 207:34]
  wire  sum_414 = sum_303 ^ sum_304; // @[Mul.scala 206:34]
  wire  cout_414 = sum_303 & sum_304; // @[Mul.scala 207:34]
  wire  sum_415 = cout_301 ^ cout_302; // @[Mul.scala 206:34]
  wire  cout_415 = cout_301 & cout_302; // @[Mul.scala 207:34]
  wire  sum_416 = sum_305 ^ sum_306; // @[Mul.scala 206:34]
  wire  cout_416 = sum_305 & sum_306; // @[Mul.scala 207:34]
  wire  sum_417 = cout_303 ^ cout_304; // @[Mul.scala 206:34]
  wire  cout_417 = cout_303 & cout_304; // @[Mul.scala 207:34]
  wire  sum_418 = sum_307 ^ sum_308; // @[Mul.scala 206:34]
  wire  cout_418 = sum_307 & sum_308; // @[Mul.scala 207:34]
  wire  sum_419 = cout_305 ^ cout_306; // @[Mul.scala 206:34]
  wire  cout_419 = cout_305 & cout_306; // @[Mul.scala 207:34]
  wire  _sum_T_1028 = sum_309 ^ cout_307; // @[Mul.scala 191:34]
  wire  sum_420 = sum_309 ^ cout_307 ^ cout_308; // @[Mul.scala 191:42]
  wire  cout_420 = sum_309 & cout_307 | _sum_T_1028 & cout_308; // @[Mul.scala 192:44]
  wire  sum_421 = sum_310 ^ cout_309; // @[Mul.scala 206:34]
  wire  cout_421 = sum_310 & cout_309; // @[Mul.scala 207:34]
  wire  sum_422 = sum_311 ^ cout_310; // @[Mul.scala 206:34]
  wire  cout_422 = sum_311 & cout_310; // @[Mul.scala 207:34]
  wire  sum_423 = sum_312 ^ cout_311; // @[Mul.scala 206:34]
  wire  cout_423 = sum_312 & cout_311; // @[Mul.scala 207:34]
  wire  sum_424 = sum_313 ^ cout_312; // @[Mul.scala 206:34]
  wire  cout_424 = sum_313 & cout_312; // @[Mul.scala 207:34]
  wire  sum_425 = sum_314 ^ cout_313; // @[Mul.scala 206:34]
  wire  sum_432 = sum_321 ^ cout_320; // @[Mul.scala 206:34]
  wire  cout_432 = sum_321 & cout_320; // @[Mul.scala 207:34]
  wire  sum_433 = sum_322 ^ cout_321; // @[Mul.scala 206:34]
  wire  cout_433 = sum_322 & cout_321; // @[Mul.scala 207:34]
  wire  sum_434 = sum_323 ^ cout_322; // @[Mul.scala 206:34]
  wire  cout_434 = sum_323 & cout_322; // @[Mul.scala 207:34]
  wire  _sum_T_1044 = sum_324 ^ sum_325; // @[Mul.scala 191:34]
  wire  sum_435 = sum_324 ^ sum_325 ^ cout_323; // @[Mul.scala 191:42]
  wire  cout_435 = sum_324 & sum_325 | _sum_T_1044 & cout_323; // @[Mul.scala 192:44]
  wire  sum_436 = sum_326 ^ sum_327; // @[Mul.scala 206:34]
  wire  cout_436 = sum_326 & sum_327; // @[Mul.scala 207:34]
  wire  sum_437 = cout_324 ^ cout_325; // @[Mul.scala 206:34]
  wire  cout_437 = cout_324 & cout_325; // @[Mul.scala 207:34]
  wire  sum_438 = sum_328 ^ sum_329; // @[Mul.scala 206:34]
  wire  cout_438 = sum_328 & sum_329; // @[Mul.scala 207:34]
  wire  sum_439 = cout_326 ^ cout_327; // @[Mul.scala 206:34]
  wire  cout_439 = cout_326 & cout_327; // @[Mul.scala 207:34]
  wire  sum_440 = sum_330 ^ sum_331; // @[Mul.scala 206:34]
  wire  cout_440 = sum_330 & sum_331; // @[Mul.scala 207:34]
  wire  sum_441 = cout_328 ^ cout_329; // @[Mul.scala 206:34]
  wire  cout_441 = cout_328 & cout_329; // @[Mul.scala 207:34]
  wire  sum_442 = sum_332 ^ sum_333; // @[Mul.scala 206:34]
  wire  cout_442 = sum_332 & sum_333; // @[Mul.scala 207:34]
  wire  sum_443 = cout_330 ^ cout_331; // @[Mul.scala 206:34]
  wire  cout_443 = cout_330 & cout_331; // @[Mul.scala 207:34]
  wire  sum_444 = sum_334 ^ sum_335; // @[Mul.scala 206:34]
  wire  cout_444 = sum_334 & sum_335; // @[Mul.scala 207:34]
  wire  sum_445 = cout_332 ^ cout_333; // @[Mul.scala 206:34]
  wire  cout_445 = cout_332 & cout_333; // @[Mul.scala 207:34]
  wire  sum_446 = sum_336 ^ sum_337; // @[Mul.scala 206:34]
  wire  cout_446 = sum_336 & sum_337; // @[Mul.scala 207:34]
  wire  sum_447 = cout_334 ^ cout_335; // @[Mul.scala 206:34]
  wire  cout_447 = cout_334 & cout_335; // @[Mul.scala 207:34]
  wire  sum_448 = sum_338 ^ sum_339; // @[Mul.scala 206:34]
  wire  cout_448 = sum_338 & sum_339; // @[Mul.scala 207:34]
  wire  sum_449 = cout_336 ^ cout_337; // @[Mul.scala 206:34]
  wire  cout_449 = cout_336 & cout_337; // @[Mul.scala 207:34]
  wire  sum_450 = sum_340 ^ sum_341; // @[Mul.scala 206:34]
  wire  cout_450 = sum_340 & sum_341; // @[Mul.scala 207:34]
  wire  sum_451 = cout_338 ^ cout_339; // @[Mul.scala 206:34]
  wire  cout_451 = cout_338 & cout_339; // @[Mul.scala 207:34]
  wire  sum_452 = sum_342 ^ sum_343; // @[Mul.scala 206:34]
  wire  cout_452 = sum_342 & sum_343; // @[Mul.scala 207:34]
  wire  sum_453 = cout_340 ^ cout_341; // @[Mul.scala 206:34]
  wire  cout_453 = cout_340 & cout_341; // @[Mul.scala 207:34]
  wire  sum_454 = sum_344 ^ sum_345; // @[Mul.scala 206:34]
  wire  cout_454 = sum_344 & sum_345; // @[Mul.scala 207:34]
  wire  sum_455 = cout_342 ^ cout_343; // @[Mul.scala 206:34]
  wire  cout_455 = cout_342 & cout_343; // @[Mul.scala 207:34]
  wire  sum_456 = sum_346 ^ sum_347; // @[Mul.scala 206:34]
  wire  cout_456 = sum_346 & sum_347; // @[Mul.scala 207:34]
  wire  sum_457 = cout_344 ^ cout_345; // @[Mul.scala 206:34]
  wire  cout_457 = cout_344 & cout_345; // @[Mul.scala 207:34]
  wire  sum_458 = sum_348 ^ sum_349; // @[Mul.scala 206:34]
  wire  cout_458 = sum_348 & sum_349; // @[Mul.scala 207:34]
  wire  sum_459 = cout_346 ^ cout_347; // @[Mul.scala 206:34]
  wire  cout_459 = cout_346 & cout_347; // @[Mul.scala 207:34]
  wire  sum_460 = sum_350 ^ sum_351; // @[Mul.scala 206:34]
  wire  cout_460 = sum_350 & sum_351; // @[Mul.scala 207:34]
  wire  sum_461 = cout_348 ^ cout_349; // @[Mul.scala 206:34]
  wire  cout_461 = cout_348 & cout_349; // @[Mul.scala 207:34]
  wire  sum_462 = sum_352 ^ sum_353; // @[Mul.scala 206:34]
  wire  cout_462 = sum_352 & sum_353; // @[Mul.scala 207:34]
  wire  sum_463 = cout_350 ^ cout_351; // @[Mul.scala 206:34]
  wire  cout_463 = cout_350 & cout_351; // @[Mul.scala 207:34]
  wire  sum_464 = sum_354 ^ sum_355; // @[Mul.scala 206:34]
  wire  cout_464 = sum_354 & sum_355; // @[Mul.scala 207:34]
  wire  sum_465 = cout_352 ^ cout_353; // @[Mul.scala 206:34]
  wire  cout_465 = cout_352 & cout_353; // @[Mul.scala 207:34]
  wire  sum_466 = sum_356 ^ sum_357; // @[Mul.scala 206:34]
  wire  cout_466 = sum_356 & sum_357; // @[Mul.scala 207:34]
  wire  sum_467 = cout_354 ^ cout_355; // @[Mul.scala 206:34]
  wire  cout_467 = cout_354 & cout_355; // @[Mul.scala 207:34]
  wire  sum_468 = sum_358 ^ sum_359; // @[Mul.scala 206:34]
  wire  cout_468 = sum_358 & sum_359; // @[Mul.scala 207:34]
  wire  sum_469 = cout_356 ^ cout_357; // @[Mul.scala 206:34]
  wire  cout_469 = cout_356 & cout_357; // @[Mul.scala 207:34]
  wire  sum_470 = sum_360 ^ sum_361; // @[Mul.scala 206:34]
  wire  cout_470 = sum_360 & sum_361; // @[Mul.scala 207:34]
  wire  sum_471 = cout_358 ^ cout_359; // @[Mul.scala 206:34]
  wire  cout_471 = cout_358 & cout_359; // @[Mul.scala 207:34]
  wire  sum_472 = sum_362 ^ sum_363; // @[Mul.scala 206:34]
  wire  cout_472 = sum_362 & sum_363; // @[Mul.scala 207:34]
  wire  sum_473 = cout_360 ^ cout_361; // @[Mul.scala 206:34]
  wire  cout_473 = cout_360 & cout_361; // @[Mul.scala 207:34]
  wire  sum_474 = sum_364 ^ sum_365; // @[Mul.scala 206:34]
  wire  cout_474 = sum_364 & sum_365; // @[Mul.scala 207:34]
  wire  sum_475 = cout_362 ^ cout_363; // @[Mul.scala 206:34]
  wire  cout_475 = cout_362 & cout_363; // @[Mul.scala 207:34]
  wire  sum_476 = sum_366 ^ sum_367; // @[Mul.scala 206:34]
  wire  cout_476 = sum_366 & sum_367; // @[Mul.scala 207:34]
  wire  sum_477 = cout_364 ^ cout_365; // @[Mul.scala 206:34]
  wire  cout_477 = cout_364 & cout_365; // @[Mul.scala 207:34]
  wire  sum_478 = sum_368 ^ sum_369; // @[Mul.scala 206:34]
  wire  cout_478 = sum_368 & sum_369; // @[Mul.scala 207:34]
  wire  sum_479 = cout_366 ^ cout_367; // @[Mul.scala 206:34]
  wire  cout_479 = cout_366 & cout_367; // @[Mul.scala 207:34]
  wire  sum_480 = sum_370 ^ sum_371; // @[Mul.scala 206:34]
  wire  cout_480 = sum_370 & sum_371; // @[Mul.scala 207:34]
  wire  sum_481 = cout_368 ^ cout_369; // @[Mul.scala 206:34]
  wire  cout_481 = cout_368 & cout_369; // @[Mul.scala 207:34]
  wire  sum_482 = sum_372 ^ sum_373; // @[Mul.scala 206:34]
  wire  cout_482 = sum_372 & sum_373; // @[Mul.scala 207:34]
  wire  sum_483 = cout_370 ^ cout_371; // @[Mul.scala 206:34]
  wire  cout_483 = cout_370 & cout_371; // @[Mul.scala 207:34]
  wire  sum_484 = sum_374 ^ sum_375; // @[Mul.scala 206:34]
  wire  cout_484 = sum_374 & sum_375; // @[Mul.scala 207:34]
  wire  sum_485 = cout_372 ^ cout_373; // @[Mul.scala 206:34]
  wire  cout_485 = cout_372 & cout_373; // @[Mul.scala 207:34]
  wire  sum_486 = sum_376 ^ sum_377; // @[Mul.scala 206:34]
  wire  cout_486 = sum_376 & sum_377; // @[Mul.scala 207:34]
  wire  sum_487 = cout_374 ^ cout_375; // @[Mul.scala 206:34]
  wire  cout_487 = cout_374 & cout_375; // @[Mul.scala 207:34]
  wire  sum_488 = sum_378 ^ sum_379; // @[Mul.scala 206:34]
  wire  cout_488 = sum_378 & sum_379; // @[Mul.scala 207:34]
  wire  sum_489 = cout_376 ^ cout_377; // @[Mul.scala 206:34]
  wire  cout_489 = cout_376 & cout_377; // @[Mul.scala 207:34]
  wire  sum_490 = sum_380 ^ sum_381; // @[Mul.scala 206:34]
  wire  cout_490 = sum_380 & sum_381; // @[Mul.scala 207:34]
  wire  sum_491 = cout_378 ^ cout_379; // @[Mul.scala 206:34]
  wire  cout_491 = cout_378 & cout_379; // @[Mul.scala 207:34]
  wire  sum_492 = sum_382 ^ sum_383; // @[Mul.scala 206:34]
  wire  cout_492 = sum_382 & sum_383; // @[Mul.scala 207:34]
  wire  sum_493 = cout_380 ^ cout_381; // @[Mul.scala 206:34]
  wire  cout_493 = cout_380 & cout_381; // @[Mul.scala 207:34]
  wire  sum_494 = sum_384 ^ sum_385; // @[Mul.scala 206:34]
  wire  cout_494 = sum_384 & sum_385; // @[Mul.scala 207:34]
  wire  sum_495 = cout_382 ^ cout_383; // @[Mul.scala 206:34]
  wire  cout_495 = cout_382 & cout_383; // @[Mul.scala 207:34]
  wire  sum_496 = sum_386 ^ sum_387; // @[Mul.scala 206:34]
  wire  cout_496 = sum_386 & sum_387; // @[Mul.scala 207:34]
  wire  sum_497 = cout_384 ^ cout_385; // @[Mul.scala 206:34]
  wire  cout_497 = cout_384 & cout_385; // @[Mul.scala 207:34]
  wire  sum_498 = sum_388 ^ sum_389; // @[Mul.scala 206:34]
  wire  cout_498 = sum_388 & sum_389; // @[Mul.scala 207:34]
  wire  sum_499 = cout_386 ^ cout_387; // @[Mul.scala 206:34]
  wire  cout_499 = cout_386 & cout_387; // @[Mul.scala 207:34]
  wire  sum_500 = sum_390 ^ sum_391; // @[Mul.scala 206:34]
  wire  cout_500 = sum_390 & sum_391; // @[Mul.scala 207:34]
  wire  sum_501 = cout_388 ^ cout_389; // @[Mul.scala 206:34]
  wire  cout_501 = cout_388 & cout_389; // @[Mul.scala 207:34]
  wire  sum_502 = sum_392 ^ sum_393; // @[Mul.scala 206:34]
  wire  cout_502 = sum_392 & sum_393; // @[Mul.scala 207:34]
  wire  sum_503 = cout_390 ^ cout_391; // @[Mul.scala 206:34]
  wire  cout_503 = cout_390 & cout_391; // @[Mul.scala 207:34]
  wire  sum_504 = sum_394 ^ sum_395; // @[Mul.scala 206:34]
  wire  cout_504 = sum_394 & sum_395; // @[Mul.scala 207:34]
  wire  sum_505 = cout_392 ^ cout_393; // @[Mul.scala 206:34]
  wire  cout_505 = cout_392 & cout_393; // @[Mul.scala 207:34]
  wire  sum_506 = sum_396 ^ sum_397; // @[Mul.scala 206:34]
  wire  cout_506 = sum_396 & sum_397; // @[Mul.scala 207:34]
  wire  sum_507 = cout_394 ^ cout_395; // @[Mul.scala 206:34]
  wire  cout_507 = cout_394 & cout_395; // @[Mul.scala 207:34]
  wire  sum_508 = sum_398 ^ sum_399; // @[Mul.scala 206:34]
  wire  cout_508 = sum_398 & sum_399; // @[Mul.scala 207:34]
  wire  sum_509 = cout_396 ^ cout_397; // @[Mul.scala 206:34]
  wire  cout_509 = cout_396 & cout_397; // @[Mul.scala 207:34]
  wire  sum_510 = sum_400 ^ sum_401; // @[Mul.scala 206:34]
  wire  cout_510 = sum_400 & sum_401; // @[Mul.scala 207:34]
  wire  sum_511 = cout_398 ^ cout_399; // @[Mul.scala 206:34]
  wire  cout_511 = cout_398 & cout_399; // @[Mul.scala 207:34]
  wire  sum_512 = sum_402 ^ sum_403; // @[Mul.scala 206:34]
  wire  cout_512 = sum_402 & sum_403; // @[Mul.scala 207:34]
  wire  sum_513 = cout_400 ^ cout_401; // @[Mul.scala 206:34]
  wire  cout_513 = cout_400 & cout_401; // @[Mul.scala 207:34]
  wire  sum_514 = sum_404 ^ sum_405; // @[Mul.scala 206:34]
  wire  cout_514 = sum_404 & sum_405; // @[Mul.scala 207:34]
  wire  sum_515 = cout_402 ^ cout_403; // @[Mul.scala 206:34]
  wire  cout_515 = cout_402 & cout_403; // @[Mul.scala 207:34]
  wire  sum_516 = sum_406 ^ sum_407; // @[Mul.scala 206:34]
  wire  cout_516 = sum_406 & sum_407; // @[Mul.scala 207:34]
  wire  sum_517 = cout_404 ^ cout_405; // @[Mul.scala 206:34]
  wire  cout_517 = cout_404 & cout_405; // @[Mul.scala 207:34]
  wire  sum_518 = sum_408 ^ sum_409; // @[Mul.scala 206:34]
  wire  cout_518 = sum_408 & sum_409; // @[Mul.scala 207:34]
  wire  sum_519 = cout_406 ^ cout_407; // @[Mul.scala 206:34]
  wire  cout_519 = cout_406 & cout_407; // @[Mul.scala 207:34]
  wire  sum_520 = sum_410 ^ sum_411; // @[Mul.scala 206:34]
  wire  cout_520 = sum_410 & sum_411; // @[Mul.scala 207:34]
  wire  sum_521 = cout_408 ^ cout_409; // @[Mul.scala 206:34]
  wire  cout_521 = cout_408 & cout_409; // @[Mul.scala 207:34]
  wire  sum_522 = sum_412 ^ sum_413; // @[Mul.scala 206:34]
  wire  cout_522 = sum_412 & sum_413; // @[Mul.scala 207:34]
  wire  sum_523 = cout_410 ^ cout_411; // @[Mul.scala 206:34]
  wire  cout_523 = cout_410 & cout_411; // @[Mul.scala 207:34]
  wire  sum_524 = sum_414 ^ sum_415; // @[Mul.scala 206:34]
  wire  cout_524 = sum_414 & sum_415; // @[Mul.scala 207:34]
  wire  sum_525 = cout_412 ^ cout_413; // @[Mul.scala 206:34]
  wire  cout_525 = cout_412 & cout_413; // @[Mul.scala 207:34]
  wire  sum_526 = sum_416 ^ sum_417; // @[Mul.scala 206:34]
  wire  cout_526 = sum_416 & sum_417; // @[Mul.scala 207:34]
  wire  sum_527 = cout_414 ^ cout_415; // @[Mul.scala 206:34]
  wire  cout_527 = cout_414 & cout_415; // @[Mul.scala 207:34]
  wire  sum_528 = sum_418 ^ sum_419; // @[Mul.scala 206:34]
  wire  cout_528 = sum_418 & sum_419; // @[Mul.scala 207:34]
  wire  sum_529 = cout_416 ^ cout_417; // @[Mul.scala 206:34]
  wire  cout_529 = cout_416 & cout_417; // @[Mul.scala 207:34]
  wire  _sum_T_1140 = sum_420 ^ cout_418; // @[Mul.scala 191:34]
  wire  sum_530 = sum_420 ^ cout_418 ^ cout_419; // @[Mul.scala 191:42]
  wire  cout_530 = sum_420 & cout_418 | _sum_T_1140 & cout_419; // @[Mul.scala 192:44]
  wire  sum_531 = sum_421 ^ cout_420; // @[Mul.scala 206:34]
  wire  cout_531 = sum_421 & cout_420; // @[Mul.scala 207:34]
  wire  sum_532 = sum_422 ^ cout_421; // @[Mul.scala 206:34]
  wire  cout_532 = sum_422 & cout_421; // @[Mul.scala 207:34]
  wire  sum_533 = sum_423 ^ cout_422; // @[Mul.scala 206:34]
  wire  cout_533 = sum_423 & cout_422; // @[Mul.scala 207:34]
  wire  sum_534 = sum_424 ^ cout_423; // @[Mul.scala 206:34]
  wire  cout_534 = sum_424 & cout_423; // @[Mul.scala 207:34]
  wire  sum_535 = sum_425 ^ cout_424; // @[Mul.scala 206:34]
  wire  sum_543 = sum_433 ^ cout_432; // @[Mul.scala 206:34]
  wire  cout_543 = sum_433 & cout_432; // @[Mul.scala 207:34]
  wire  sum_544 = sum_434 ^ cout_433; // @[Mul.scala 206:34]
  wire  cout_544 = sum_434 & cout_433; // @[Mul.scala 207:34]
  wire  sum_545 = sum_435 ^ cout_434; // @[Mul.scala 206:34]
  wire  cout_545 = sum_435 & cout_434; // @[Mul.scala 207:34]
  wire  _sum_T_1157 = sum_436 ^ sum_437; // @[Mul.scala 191:34]
  wire  sum_546 = sum_436 ^ sum_437 ^ cout_435; // @[Mul.scala 191:42]
  wire  cout_546 = sum_436 & sum_437 | _sum_T_1157 & cout_435; // @[Mul.scala 192:44]
  wire  sum_547 = sum_438 ^ sum_439; // @[Mul.scala 206:34]
  wire  cout_547 = sum_438 & sum_439; // @[Mul.scala 207:34]
  wire  sum_548 = cout_436 ^ cout_437; // @[Mul.scala 206:34]
  wire  cout_548 = cout_436 & cout_437; // @[Mul.scala 207:34]
  wire  sum_549 = sum_440 ^ sum_441; // @[Mul.scala 206:34]
  wire  cout_549 = sum_440 & sum_441; // @[Mul.scala 207:34]
  wire  sum_550 = cout_438 ^ cout_439; // @[Mul.scala 206:34]
  wire  cout_550 = cout_438 & cout_439; // @[Mul.scala 207:34]
  wire  sum_551 = sum_442 ^ sum_443; // @[Mul.scala 206:34]
  wire  cout_551 = sum_442 & sum_443; // @[Mul.scala 207:34]
  wire  sum_552 = cout_440 ^ cout_441; // @[Mul.scala 206:34]
  wire  cout_552 = cout_440 & cout_441; // @[Mul.scala 207:34]
  wire  sum_553 = sum_444 ^ sum_445; // @[Mul.scala 206:34]
  wire  cout_553 = sum_444 & sum_445; // @[Mul.scala 207:34]
  wire  sum_554 = cout_442 ^ cout_443; // @[Mul.scala 206:34]
  wire  cout_554 = cout_442 & cout_443; // @[Mul.scala 207:34]
  wire  sum_555 = sum_446 ^ sum_447; // @[Mul.scala 206:34]
  wire  cout_555 = sum_446 & sum_447; // @[Mul.scala 207:34]
  wire  sum_556 = cout_444 ^ cout_445; // @[Mul.scala 206:34]
  wire  cout_556 = cout_444 & cout_445; // @[Mul.scala 207:34]
  wire  sum_557 = sum_448 ^ sum_449; // @[Mul.scala 206:34]
  wire  cout_557 = sum_448 & sum_449; // @[Mul.scala 207:34]
  wire  sum_558 = cout_446 ^ cout_447; // @[Mul.scala 206:34]
  wire  cout_558 = cout_446 & cout_447; // @[Mul.scala 207:34]
  wire  sum_559 = sum_450 ^ sum_451; // @[Mul.scala 206:34]
  wire  cout_559 = sum_450 & sum_451; // @[Mul.scala 207:34]
  wire  sum_560 = cout_448 ^ cout_449; // @[Mul.scala 206:34]
  wire  cout_560 = cout_448 & cout_449; // @[Mul.scala 207:34]
  wire  sum_561 = sum_452 ^ sum_453; // @[Mul.scala 206:34]
  wire  cout_561 = sum_452 & sum_453; // @[Mul.scala 207:34]
  wire  sum_562 = cout_450 ^ cout_451; // @[Mul.scala 206:34]
  wire  cout_562 = cout_450 & cout_451; // @[Mul.scala 207:34]
  wire  sum_563 = sum_454 ^ sum_455; // @[Mul.scala 206:34]
  wire  cout_563 = sum_454 & sum_455; // @[Mul.scala 207:34]
  wire  sum_564 = cout_452 ^ cout_453; // @[Mul.scala 206:34]
  wire  cout_564 = cout_452 & cout_453; // @[Mul.scala 207:34]
  wire  sum_565 = sum_456 ^ sum_457; // @[Mul.scala 206:34]
  wire  cout_565 = sum_456 & sum_457; // @[Mul.scala 207:34]
  wire  sum_566 = cout_454 ^ cout_455; // @[Mul.scala 206:34]
  wire  cout_566 = cout_454 & cout_455; // @[Mul.scala 207:34]
  wire  sum_567 = sum_458 ^ sum_459; // @[Mul.scala 206:34]
  wire  cout_567 = sum_458 & sum_459; // @[Mul.scala 207:34]
  wire  sum_568 = cout_456 ^ cout_457; // @[Mul.scala 206:34]
  wire  cout_568 = cout_456 & cout_457; // @[Mul.scala 207:34]
  wire  sum_569 = sum_460 ^ sum_461; // @[Mul.scala 206:34]
  wire  cout_569 = sum_460 & sum_461; // @[Mul.scala 207:34]
  wire  sum_570 = cout_458 ^ cout_459; // @[Mul.scala 206:34]
  wire  cout_570 = cout_458 & cout_459; // @[Mul.scala 207:34]
  wire  sum_571 = sum_462 ^ sum_463; // @[Mul.scala 206:34]
  wire  cout_571 = sum_462 & sum_463; // @[Mul.scala 207:34]
  wire  sum_572 = cout_460 ^ cout_461; // @[Mul.scala 206:34]
  wire  cout_572 = cout_460 & cout_461; // @[Mul.scala 207:34]
  wire  sum_573 = sum_464 ^ sum_465; // @[Mul.scala 206:34]
  wire  cout_573 = sum_464 & sum_465; // @[Mul.scala 207:34]
  wire  sum_574 = cout_462 ^ cout_463; // @[Mul.scala 206:34]
  wire  cout_574 = cout_462 & cout_463; // @[Mul.scala 207:34]
  wire  sum_575 = sum_466 ^ sum_467; // @[Mul.scala 206:34]
  wire  cout_575 = sum_466 & sum_467; // @[Mul.scala 207:34]
  wire  sum_576 = cout_464 ^ cout_465; // @[Mul.scala 206:34]
  wire  cout_576 = cout_464 & cout_465; // @[Mul.scala 207:34]
  wire  sum_577 = sum_468 ^ sum_469; // @[Mul.scala 206:34]
  wire  cout_577 = sum_468 & sum_469; // @[Mul.scala 207:34]
  wire  sum_578 = cout_466 ^ cout_467; // @[Mul.scala 206:34]
  wire  cout_578 = cout_466 & cout_467; // @[Mul.scala 207:34]
  wire  sum_579 = sum_470 ^ sum_471; // @[Mul.scala 206:34]
  wire  cout_579 = sum_470 & sum_471; // @[Mul.scala 207:34]
  wire  sum_580 = cout_468 ^ cout_469; // @[Mul.scala 206:34]
  wire  cout_580 = cout_468 & cout_469; // @[Mul.scala 207:34]
  wire  sum_581 = sum_472 ^ sum_473; // @[Mul.scala 206:34]
  wire  cout_581 = sum_472 & sum_473; // @[Mul.scala 207:34]
  wire  sum_582 = cout_470 ^ cout_471; // @[Mul.scala 206:34]
  wire  cout_582 = cout_470 & cout_471; // @[Mul.scala 207:34]
  wire  sum_583 = sum_474 ^ sum_475; // @[Mul.scala 206:34]
  wire  cout_583 = sum_474 & sum_475; // @[Mul.scala 207:34]
  wire  sum_584 = cout_472 ^ cout_473; // @[Mul.scala 206:34]
  wire  cout_584 = cout_472 & cout_473; // @[Mul.scala 207:34]
  wire  sum_585 = sum_476 ^ sum_477; // @[Mul.scala 206:34]
  wire  cout_585 = sum_476 & sum_477; // @[Mul.scala 207:34]
  wire  sum_586 = cout_474 ^ cout_475; // @[Mul.scala 206:34]
  wire  cout_586 = cout_474 & cout_475; // @[Mul.scala 207:34]
  wire  sum_587 = sum_478 ^ sum_479; // @[Mul.scala 206:34]
  wire  cout_587 = sum_478 & sum_479; // @[Mul.scala 207:34]
  wire  sum_588 = cout_476 ^ cout_477; // @[Mul.scala 206:34]
  wire  cout_588 = cout_476 & cout_477; // @[Mul.scala 207:34]
  wire  sum_589 = sum_480 ^ sum_481; // @[Mul.scala 206:34]
  wire  cout_589 = sum_480 & sum_481; // @[Mul.scala 207:34]
  wire  sum_590 = cout_478 ^ cout_479; // @[Mul.scala 206:34]
  wire  cout_590 = cout_478 & cout_479; // @[Mul.scala 207:34]
  wire  sum_591 = sum_482 ^ sum_483; // @[Mul.scala 206:34]
  wire  cout_591 = sum_482 & sum_483; // @[Mul.scala 207:34]
  wire  sum_592 = cout_480 ^ cout_481; // @[Mul.scala 206:34]
  wire  cout_592 = cout_480 & cout_481; // @[Mul.scala 207:34]
  wire  sum_593 = sum_484 ^ sum_485; // @[Mul.scala 206:34]
  wire  cout_593 = sum_484 & sum_485; // @[Mul.scala 207:34]
  wire  sum_594 = cout_482 ^ cout_483; // @[Mul.scala 206:34]
  wire  cout_594 = cout_482 & cout_483; // @[Mul.scala 207:34]
  wire  sum_595 = sum_486 ^ sum_487; // @[Mul.scala 206:34]
  wire  cout_595 = sum_486 & sum_487; // @[Mul.scala 207:34]
  wire  sum_596 = cout_484 ^ cout_485; // @[Mul.scala 206:34]
  wire  cout_596 = cout_484 & cout_485; // @[Mul.scala 207:34]
  wire  sum_597 = sum_488 ^ sum_489; // @[Mul.scala 206:34]
  wire  cout_597 = sum_488 & sum_489; // @[Mul.scala 207:34]
  wire  sum_598 = cout_486 ^ cout_487; // @[Mul.scala 206:34]
  wire  cout_598 = cout_486 & cout_487; // @[Mul.scala 207:34]
  wire  sum_599 = sum_490 ^ sum_491; // @[Mul.scala 206:34]
  wire  cout_599 = sum_490 & sum_491; // @[Mul.scala 207:34]
  wire  sum_600 = cout_488 ^ cout_489; // @[Mul.scala 206:34]
  wire  cout_600 = cout_488 & cout_489; // @[Mul.scala 207:34]
  wire  sum_601 = sum_492 ^ sum_493; // @[Mul.scala 206:34]
  wire  cout_601 = sum_492 & sum_493; // @[Mul.scala 207:34]
  wire  sum_602 = cout_490 ^ cout_491; // @[Mul.scala 206:34]
  wire  cout_602 = cout_490 & cout_491; // @[Mul.scala 207:34]
  wire  sum_603 = sum_494 ^ sum_495; // @[Mul.scala 206:34]
  wire  cout_603 = sum_494 & sum_495; // @[Mul.scala 207:34]
  wire  sum_604 = cout_492 ^ cout_493; // @[Mul.scala 206:34]
  wire  cout_604 = cout_492 & cout_493; // @[Mul.scala 207:34]
  wire  sum_605 = sum_496 ^ sum_497; // @[Mul.scala 206:34]
  wire  cout_605 = sum_496 & sum_497; // @[Mul.scala 207:34]
  wire  sum_606 = cout_494 ^ cout_495; // @[Mul.scala 206:34]
  wire  cout_606 = cout_494 & cout_495; // @[Mul.scala 207:34]
  wire  sum_607 = sum_498 ^ sum_499; // @[Mul.scala 206:34]
  wire  cout_607 = sum_498 & sum_499; // @[Mul.scala 207:34]
  wire  sum_608 = cout_496 ^ cout_497; // @[Mul.scala 206:34]
  wire  cout_608 = cout_496 & cout_497; // @[Mul.scala 207:34]
  wire  sum_609 = sum_500 ^ sum_501; // @[Mul.scala 206:34]
  wire  cout_609 = sum_500 & sum_501; // @[Mul.scala 207:34]
  wire  sum_610 = cout_498 ^ cout_499; // @[Mul.scala 206:34]
  wire  cout_610 = cout_498 & cout_499; // @[Mul.scala 207:34]
  wire  sum_611 = sum_502 ^ sum_503; // @[Mul.scala 206:34]
  wire  cout_611 = sum_502 & sum_503; // @[Mul.scala 207:34]
  wire  sum_612 = cout_500 ^ cout_501; // @[Mul.scala 206:34]
  wire  cout_612 = cout_500 & cout_501; // @[Mul.scala 207:34]
  wire  sum_613 = sum_504 ^ sum_505; // @[Mul.scala 206:34]
  wire  cout_613 = sum_504 & sum_505; // @[Mul.scala 207:34]
  wire  sum_614 = cout_502 ^ cout_503; // @[Mul.scala 206:34]
  wire  cout_614 = cout_502 & cout_503; // @[Mul.scala 207:34]
  wire  sum_615 = sum_506 ^ sum_507; // @[Mul.scala 206:34]
  wire  cout_615 = sum_506 & sum_507; // @[Mul.scala 207:34]
  wire  sum_616 = cout_504 ^ cout_505; // @[Mul.scala 206:34]
  wire  cout_616 = cout_504 & cout_505; // @[Mul.scala 207:34]
  wire  sum_617 = sum_508 ^ sum_509; // @[Mul.scala 206:34]
  wire  cout_617 = sum_508 & sum_509; // @[Mul.scala 207:34]
  wire  sum_618 = cout_506 ^ cout_507; // @[Mul.scala 206:34]
  wire  cout_618 = cout_506 & cout_507; // @[Mul.scala 207:34]
  wire  sum_619 = sum_510 ^ sum_511; // @[Mul.scala 206:34]
  wire  cout_619 = sum_510 & sum_511; // @[Mul.scala 207:34]
  wire  sum_620 = cout_508 ^ cout_509; // @[Mul.scala 206:34]
  wire  cout_620 = cout_508 & cout_509; // @[Mul.scala 207:34]
  wire  sum_621 = sum_512 ^ sum_513; // @[Mul.scala 206:34]
  wire  cout_621 = sum_512 & sum_513; // @[Mul.scala 207:34]
  wire  sum_622 = cout_510 ^ cout_511; // @[Mul.scala 206:34]
  wire  cout_622 = cout_510 & cout_511; // @[Mul.scala 207:34]
  wire  sum_623 = sum_514 ^ sum_515; // @[Mul.scala 206:34]
  wire  cout_623 = sum_514 & sum_515; // @[Mul.scala 207:34]
  wire  sum_624 = cout_512 ^ cout_513; // @[Mul.scala 206:34]
  wire  cout_624 = cout_512 & cout_513; // @[Mul.scala 207:34]
  wire  sum_625 = sum_516 ^ sum_517; // @[Mul.scala 206:34]
  wire  cout_625 = sum_516 & sum_517; // @[Mul.scala 207:34]
  wire  sum_626 = cout_514 ^ cout_515; // @[Mul.scala 206:34]
  wire  cout_626 = cout_514 & cout_515; // @[Mul.scala 207:34]
  wire  sum_627 = sum_518 ^ sum_519; // @[Mul.scala 206:34]
  wire  cout_627 = sum_518 & sum_519; // @[Mul.scala 207:34]
  wire  sum_628 = cout_516 ^ cout_517; // @[Mul.scala 206:34]
  wire  cout_628 = cout_516 & cout_517; // @[Mul.scala 207:34]
  wire  sum_629 = sum_520 ^ sum_521; // @[Mul.scala 206:34]
  wire  cout_629 = sum_520 & sum_521; // @[Mul.scala 207:34]
  wire  sum_630 = cout_518 ^ cout_519; // @[Mul.scala 206:34]
  wire  cout_630 = cout_518 & cout_519; // @[Mul.scala 207:34]
  wire  sum_631 = sum_522 ^ sum_523; // @[Mul.scala 206:34]
  wire  cout_631 = sum_522 & sum_523; // @[Mul.scala 207:34]
  wire  sum_632 = cout_520 ^ cout_521; // @[Mul.scala 206:34]
  wire  cout_632 = cout_520 & cout_521; // @[Mul.scala 207:34]
  wire  sum_633 = sum_524 ^ sum_525; // @[Mul.scala 206:34]
  wire  cout_633 = sum_524 & sum_525; // @[Mul.scala 207:34]
  wire  sum_634 = cout_522 ^ cout_523; // @[Mul.scala 206:34]
  wire  cout_634 = cout_522 & cout_523; // @[Mul.scala 207:34]
  wire  sum_635 = sum_526 ^ sum_527; // @[Mul.scala 206:34]
  wire  cout_635 = sum_526 & sum_527; // @[Mul.scala 207:34]
  wire  sum_636 = cout_524 ^ cout_525; // @[Mul.scala 206:34]
  wire  cout_636 = cout_524 & cout_525; // @[Mul.scala 207:34]
  wire  sum_637 = sum_528 ^ sum_529; // @[Mul.scala 206:34]
  wire  cout_637 = sum_528 & sum_529; // @[Mul.scala 207:34]
  wire  sum_638 = cout_526 ^ cout_527; // @[Mul.scala 206:34]
  wire  cout_638 = cout_526 & cout_527; // @[Mul.scala 207:34]
  wire  _sum_T_1251 = sum_530 ^ cout_528; // @[Mul.scala 191:34]
  wire  sum_639 = sum_530 ^ cout_528 ^ cout_529; // @[Mul.scala 191:42]
  wire  cout_639 = sum_530 & cout_528 | _sum_T_1251 & cout_529; // @[Mul.scala 192:44]
  wire  sum_640 = sum_531 ^ cout_530; // @[Mul.scala 206:34]
  wire  cout_640 = sum_531 & cout_530; // @[Mul.scala 207:34]
  wire  sum_641 = sum_532 ^ cout_531; // @[Mul.scala 206:34]
  wire  cout_641 = sum_532 & cout_531; // @[Mul.scala 207:34]
  wire  sum_642 = sum_533 ^ cout_532; // @[Mul.scala 206:34]
  wire  cout_642 = sum_533 & cout_532; // @[Mul.scala 207:34]
  wire  sum_643 = sum_534 ^ cout_533; // @[Mul.scala 206:34]
  wire  cout_643 = sum_534 & cout_533; // @[Mul.scala 207:34]
  wire  sum_644 = sum_535 ^ cout_534; // @[Mul.scala 206:34]
  wire  sum_653 = sum_544 ^ cout_543; // @[Mul.scala 206:34]
  wire  cout_653 = sum_544 & cout_543; // @[Mul.scala 207:34]
  wire  sum_654 = sum_545 ^ cout_544; // @[Mul.scala 206:34]
  wire  cout_654 = sum_545 & cout_544; // @[Mul.scala 207:34]
  wire  sum_655 = sum_546 ^ cout_545; // @[Mul.scala 206:34]
  wire  cout_655 = sum_546 & cout_545; // @[Mul.scala 207:34]
  wire  _sum_T_1269 = sum_547 ^ sum_548; // @[Mul.scala 191:34]
  wire  sum_656 = sum_547 ^ sum_548 ^ cout_546; // @[Mul.scala 191:42]
  wire  cout_656 = sum_547 & sum_548 | _sum_T_1269 & cout_546; // @[Mul.scala 192:44]
  wire  sum_657 = sum_549 ^ sum_550; // @[Mul.scala 206:34]
  wire  cout_657 = sum_549 & sum_550; // @[Mul.scala 207:34]
  wire  sum_658 = cout_547 ^ cout_548; // @[Mul.scala 206:34]
  wire  cout_658 = cout_547 & cout_548; // @[Mul.scala 207:34]
  wire  sum_659 = sum_551 ^ sum_552; // @[Mul.scala 206:34]
  wire  cout_659 = sum_551 & sum_552; // @[Mul.scala 207:34]
  wire  sum_660 = cout_549 ^ cout_550; // @[Mul.scala 206:34]
  wire  cout_660 = cout_549 & cout_550; // @[Mul.scala 207:34]
  wire  sum_661 = sum_553 ^ sum_554; // @[Mul.scala 206:34]
  wire  cout_661 = sum_553 & sum_554; // @[Mul.scala 207:34]
  wire  sum_662 = cout_551 ^ cout_552; // @[Mul.scala 206:34]
  wire  cout_662 = cout_551 & cout_552; // @[Mul.scala 207:34]
  wire  sum_663 = sum_555 ^ sum_556; // @[Mul.scala 206:34]
  wire  cout_663 = sum_555 & sum_556; // @[Mul.scala 207:34]
  wire  sum_664 = cout_553 ^ cout_554; // @[Mul.scala 206:34]
  wire  cout_664 = cout_553 & cout_554; // @[Mul.scala 207:34]
  wire  sum_665 = sum_557 ^ sum_558; // @[Mul.scala 206:34]
  wire  cout_665 = sum_557 & sum_558; // @[Mul.scala 207:34]
  wire  sum_666 = cout_555 ^ cout_556; // @[Mul.scala 206:34]
  wire  cout_666 = cout_555 & cout_556; // @[Mul.scala 207:34]
  wire  sum_667 = sum_559 ^ sum_560; // @[Mul.scala 206:34]
  wire  cout_667 = sum_559 & sum_560; // @[Mul.scala 207:34]
  wire  sum_668 = cout_557 ^ cout_558; // @[Mul.scala 206:34]
  wire  cout_668 = cout_557 & cout_558; // @[Mul.scala 207:34]
  wire  sum_669 = sum_561 ^ sum_562; // @[Mul.scala 206:34]
  wire  cout_669 = sum_561 & sum_562; // @[Mul.scala 207:34]
  wire  sum_670 = cout_559 ^ cout_560; // @[Mul.scala 206:34]
  wire  cout_670 = cout_559 & cout_560; // @[Mul.scala 207:34]
  wire  sum_671 = sum_563 ^ sum_564; // @[Mul.scala 206:34]
  wire  cout_671 = sum_563 & sum_564; // @[Mul.scala 207:34]
  wire  sum_672 = cout_561 ^ cout_562; // @[Mul.scala 206:34]
  wire  cout_672 = cout_561 & cout_562; // @[Mul.scala 207:34]
  wire  sum_673 = sum_565 ^ sum_566; // @[Mul.scala 206:34]
  wire  cout_673 = sum_565 & sum_566; // @[Mul.scala 207:34]
  wire  sum_674 = cout_563 ^ cout_564; // @[Mul.scala 206:34]
  wire  cout_674 = cout_563 & cout_564; // @[Mul.scala 207:34]
  wire  sum_675 = sum_567 ^ sum_568; // @[Mul.scala 206:34]
  wire  cout_675 = sum_567 & sum_568; // @[Mul.scala 207:34]
  wire  sum_676 = cout_565 ^ cout_566; // @[Mul.scala 206:34]
  wire  cout_676 = cout_565 & cout_566; // @[Mul.scala 207:34]
  wire  sum_677 = sum_569 ^ sum_570; // @[Mul.scala 206:34]
  wire  cout_677 = sum_569 & sum_570; // @[Mul.scala 207:34]
  wire  sum_678 = cout_567 ^ cout_568; // @[Mul.scala 206:34]
  wire  cout_678 = cout_567 & cout_568; // @[Mul.scala 207:34]
  wire  sum_679 = sum_571 ^ sum_572; // @[Mul.scala 206:34]
  wire  cout_679 = sum_571 & sum_572; // @[Mul.scala 207:34]
  wire  sum_680 = cout_569 ^ cout_570; // @[Mul.scala 206:34]
  wire  cout_680 = cout_569 & cout_570; // @[Mul.scala 207:34]
  wire  sum_681 = sum_573 ^ sum_574; // @[Mul.scala 206:34]
  wire  cout_681 = sum_573 & sum_574; // @[Mul.scala 207:34]
  wire  sum_682 = cout_571 ^ cout_572; // @[Mul.scala 206:34]
  wire  cout_682 = cout_571 & cout_572; // @[Mul.scala 207:34]
  wire  sum_683 = sum_575 ^ sum_576; // @[Mul.scala 206:34]
  wire  cout_683 = sum_575 & sum_576; // @[Mul.scala 207:34]
  wire  sum_684 = cout_573 ^ cout_574; // @[Mul.scala 206:34]
  wire  cout_684 = cout_573 & cout_574; // @[Mul.scala 207:34]
  wire  sum_685 = sum_577 ^ sum_578; // @[Mul.scala 206:34]
  wire  cout_685 = sum_577 & sum_578; // @[Mul.scala 207:34]
  wire  sum_686 = cout_575 ^ cout_576; // @[Mul.scala 206:34]
  wire  cout_686 = cout_575 & cout_576; // @[Mul.scala 207:34]
  wire  sum_687 = sum_579 ^ sum_580; // @[Mul.scala 206:34]
  wire  cout_687 = sum_579 & sum_580; // @[Mul.scala 207:34]
  wire  sum_688 = cout_577 ^ cout_578; // @[Mul.scala 206:34]
  wire  cout_688 = cout_577 & cout_578; // @[Mul.scala 207:34]
  wire  sum_689 = sum_581 ^ sum_582; // @[Mul.scala 206:34]
  wire  cout_689 = sum_581 & sum_582; // @[Mul.scala 207:34]
  wire  sum_690 = cout_579 ^ cout_580; // @[Mul.scala 206:34]
  wire  cout_690 = cout_579 & cout_580; // @[Mul.scala 207:34]
  wire  sum_691 = sum_583 ^ sum_584; // @[Mul.scala 206:34]
  wire  cout_691 = sum_583 & sum_584; // @[Mul.scala 207:34]
  wire  sum_692 = cout_581 ^ cout_582; // @[Mul.scala 206:34]
  wire  cout_692 = cout_581 & cout_582; // @[Mul.scala 207:34]
  wire  sum_693 = sum_585 ^ sum_586; // @[Mul.scala 206:34]
  wire  cout_693 = sum_585 & sum_586; // @[Mul.scala 207:34]
  wire  sum_694 = cout_583 ^ cout_584; // @[Mul.scala 206:34]
  wire  cout_694 = cout_583 & cout_584; // @[Mul.scala 207:34]
  wire  sum_695 = sum_587 ^ sum_588; // @[Mul.scala 206:34]
  wire  cout_695 = sum_587 & sum_588; // @[Mul.scala 207:34]
  wire  sum_696 = cout_585 ^ cout_586; // @[Mul.scala 206:34]
  wire  cout_696 = cout_585 & cout_586; // @[Mul.scala 207:34]
  wire  sum_697 = sum_589 ^ sum_590; // @[Mul.scala 206:34]
  wire  cout_697 = sum_589 & sum_590; // @[Mul.scala 207:34]
  wire  sum_698 = cout_587 ^ cout_588; // @[Mul.scala 206:34]
  wire  cout_698 = cout_587 & cout_588; // @[Mul.scala 207:34]
  wire  sum_699 = sum_591 ^ sum_592; // @[Mul.scala 206:34]
  wire  cout_699 = sum_591 & sum_592; // @[Mul.scala 207:34]
  wire  sum_700 = cout_589 ^ cout_590; // @[Mul.scala 206:34]
  wire  cout_700 = cout_589 & cout_590; // @[Mul.scala 207:34]
  wire  sum_701 = sum_593 ^ sum_594; // @[Mul.scala 206:34]
  wire  cout_701 = sum_593 & sum_594; // @[Mul.scala 207:34]
  wire  sum_702 = cout_591 ^ cout_592; // @[Mul.scala 206:34]
  wire  cout_702 = cout_591 & cout_592; // @[Mul.scala 207:34]
  wire  sum_703 = sum_595 ^ sum_596; // @[Mul.scala 206:34]
  wire  cout_703 = sum_595 & sum_596; // @[Mul.scala 207:34]
  wire  sum_704 = cout_593 ^ cout_594; // @[Mul.scala 206:34]
  wire  cout_704 = cout_593 & cout_594; // @[Mul.scala 207:34]
  wire  sum_705 = sum_597 ^ sum_598; // @[Mul.scala 206:34]
  wire  cout_705 = sum_597 & sum_598; // @[Mul.scala 207:34]
  wire  sum_706 = cout_595 ^ cout_596; // @[Mul.scala 206:34]
  wire  cout_706 = cout_595 & cout_596; // @[Mul.scala 207:34]
  wire  sum_707 = sum_599 ^ sum_600; // @[Mul.scala 206:34]
  wire  cout_707 = sum_599 & sum_600; // @[Mul.scala 207:34]
  wire  sum_708 = cout_597 ^ cout_598; // @[Mul.scala 206:34]
  wire  cout_708 = cout_597 & cout_598; // @[Mul.scala 207:34]
  wire  sum_709 = sum_601 ^ sum_602; // @[Mul.scala 206:34]
  wire  cout_709 = sum_601 & sum_602; // @[Mul.scala 207:34]
  wire  sum_710 = cout_599 ^ cout_600; // @[Mul.scala 206:34]
  wire  cout_710 = cout_599 & cout_600; // @[Mul.scala 207:34]
  wire  sum_711 = sum_603 ^ sum_604; // @[Mul.scala 206:34]
  wire  cout_711 = sum_603 & sum_604; // @[Mul.scala 207:34]
  wire  sum_712 = cout_601 ^ cout_602; // @[Mul.scala 206:34]
  wire  cout_712 = cout_601 & cout_602; // @[Mul.scala 207:34]
  wire  sum_713 = sum_605 ^ sum_606; // @[Mul.scala 206:34]
  wire  cout_713 = sum_605 & sum_606; // @[Mul.scala 207:34]
  wire  sum_714 = cout_603 ^ cout_604; // @[Mul.scala 206:34]
  wire  cout_714 = cout_603 & cout_604; // @[Mul.scala 207:34]
  wire  sum_715 = sum_607 ^ sum_608; // @[Mul.scala 206:34]
  wire  cout_715 = sum_607 & sum_608; // @[Mul.scala 207:34]
  wire  sum_716 = cout_605 ^ cout_606; // @[Mul.scala 206:34]
  wire  cout_716 = cout_605 & cout_606; // @[Mul.scala 207:34]
  wire  sum_717 = sum_609 ^ sum_610; // @[Mul.scala 206:34]
  wire  cout_717 = sum_609 & sum_610; // @[Mul.scala 207:34]
  wire  sum_718 = cout_607 ^ cout_608; // @[Mul.scala 206:34]
  wire  cout_718 = cout_607 & cout_608; // @[Mul.scala 207:34]
  wire  sum_719 = sum_611 ^ sum_612; // @[Mul.scala 206:34]
  wire  cout_719 = sum_611 & sum_612; // @[Mul.scala 207:34]
  wire  sum_720 = cout_609 ^ cout_610; // @[Mul.scala 206:34]
  wire  cout_720 = cout_609 & cout_610; // @[Mul.scala 207:34]
  wire  sum_721 = sum_613 ^ sum_614; // @[Mul.scala 206:34]
  wire  cout_721 = sum_613 & sum_614; // @[Mul.scala 207:34]
  wire  sum_722 = cout_611 ^ cout_612; // @[Mul.scala 206:34]
  wire  cout_722 = cout_611 & cout_612; // @[Mul.scala 207:34]
  wire  sum_723 = sum_615 ^ sum_616; // @[Mul.scala 206:34]
  wire  cout_723 = sum_615 & sum_616; // @[Mul.scala 207:34]
  wire  sum_724 = cout_613 ^ cout_614; // @[Mul.scala 206:34]
  wire  cout_724 = cout_613 & cout_614; // @[Mul.scala 207:34]
  wire  sum_725 = sum_617 ^ sum_618; // @[Mul.scala 206:34]
  wire  cout_725 = sum_617 & sum_618; // @[Mul.scala 207:34]
  wire  sum_726 = cout_615 ^ cout_616; // @[Mul.scala 206:34]
  wire  cout_726 = cout_615 & cout_616; // @[Mul.scala 207:34]
  wire  sum_727 = sum_619 ^ sum_620; // @[Mul.scala 206:34]
  wire  cout_727 = sum_619 & sum_620; // @[Mul.scala 207:34]
  wire  sum_728 = cout_617 ^ cout_618; // @[Mul.scala 206:34]
  wire  cout_728 = cout_617 & cout_618; // @[Mul.scala 207:34]
  wire  sum_729 = sum_621 ^ sum_622; // @[Mul.scala 206:34]
  wire  cout_729 = sum_621 & sum_622; // @[Mul.scala 207:34]
  wire  sum_730 = cout_619 ^ cout_620; // @[Mul.scala 206:34]
  wire  cout_730 = cout_619 & cout_620; // @[Mul.scala 207:34]
  wire  sum_731 = sum_623 ^ sum_624; // @[Mul.scala 206:34]
  wire  cout_731 = sum_623 & sum_624; // @[Mul.scala 207:34]
  wire  sum_732 = cout_621 ^ cout_622; // @[Mul.scala 206:34]
  wire  cout_732 = cout_621 & cout_622; // @[Mul.scala 207:34]
  wire  sum_733 = sum_625 ^ sum_626; // @[Mul.scala 206:34]
  wire  cout_733 = sum_625 & sum_626; // @[Mul.scala 207:34]
  wire  sum_734 = cout_623 ^ cout_624; // @[Mul.scala 206:34]
  wire  cout_734 = cout_623 & cout_624; // @[Mul.scala 207:34]
  wire  sum_735 = sum_627 ^ sum_628; // @[Mul.scala 206:34]
  wire  cout_735 = sum_627 & sum_628; // @[Mul.scala 207:34]
  wire  sum_736 = cout_625 ^ cout_626; // @[Mul.scala 206:34]
  wire  cout_736 = cout_625 & cout_626; // @[Mul.scala 207:34]
  wire  sum_737 = sum_629 ^ sum_630; // @[Mul.scala 206:34]
  wire  cout_737 = sum_629 & sum_630; // @[Mul.scala 207:34]
  wire  sum_738 = cout_627 ^ cout_628; // @[Mul.scala 206:34]
  wire  cout_738 = cout_627 & cout_628; // @[Mul.scala 207:34]
  wire  sum_739 = sum_631 ^ sum_632; // @[Mul.scala 206:34]
  wire  cout_739 = sum_631 & sum_632; // @[Mul.scala 207:34]
  wire  sum_740 = cout_629 ^ cout_630; // @[Mul.scala 206:34]
  wire  cout_740 = cout_629 & cout_630; // @[Mul.scala 207:34]
  wire  sum_741 = sum_633 ^ sum_634; // @[Mul.scala 206:34]
  wire  cout_741 = sum_633 & sum_634; // @[Mul.scala 207:34]
  wire  sum_742 = cout_631 ^ cout_632; // @[Mul.scala 206:34]
  wire  cout_742 = cout_631 & cout_632; // @[Mul.scala 207:34]
  wire  sum_743 = sum_635 ^ sum_636; // @[Mul.scala 206:34]
  wire  cout_743 = sum_635 & sum_636; // @[Mul.scala 207:34]
  wire  sum_744 = cout_633 ^ cout_634; // @[Mul.scala 206:34]
  wire  cout_744 = cout_633 & cout_634; // @[Mul.scala 207:34]
  wire  sum_745 = sum_637 ^ sum_638; // @[Mul.scala 206:34]
  wire  cout_745 = sum_637 & sum_638; // @[Mul.scala 207:34]
  wire  sum_746 = cout_635 ^ cout_636; // @[Mul.scala 206:34]
  wire  cout_746 = cout_635 & cout_636; // @[Mul.scala 207:34]
  wire  _sum_T_1361 = sum_639 ^ cout_637; // @[Mul.scala 191:34]
  wire  sum_747 = sum_639 ^ cout_637 ^ cout_638; // @[Mul.scala 191:42]
  wire  cout_747 = sum_639 & cout_637 | _sum_T_1361 & cout_638; // @[Mul.scala 192:44]
  wire  sum_748 = sum_640 ^ cout_639; // @[Mul.scala 206:34]
  wire  cout_748 = sum_640 & cout_639; // @[Mul.scala 207:34]
  wire  sum_749 = sum_641 ^ cout_640; // @[Mul.scala 206:34]
  wire  cout_749 = sum_641 & cout_640; // @[Mul.scala 207:34]
  wire  sum_750 = sum_642 ^ cout_641; // @[Mul.scala 206:34]
  wire  cout_750 = sum_642 & cout_641; // @[Mul.scala 207:34]
  wire  sum_751 = sum_643 ^ cout_642; // @[Mul.scala 206:34]
  wire  cout_751 = sum_643 & cout_642; // @[Mul.scala 207:34]
  wire  sum_752 = sum_644 ^ cout_643; // @[Mul.scala 206:34]
  wire  sum_762 = sum_654 ^ cout_653; // @[Mul.scala 206:34]
  wire  cout_762 = sum_654 & cout_653; // @[Mul.scala 207:34]
  wire  sum_763 = sum_655 ^ cout_654; // @[Mul.scala 206:34]
  wire  cout_763 = sum_655 & cout_654; // @[Mul.scala 207:34]
  wire  sum_764 = sum_656 ^ cout_655; // @[Mul.scala 206:34]
  wire  cout_764 = sum_656 & cout_655; // @[Mul.scala 207:34]
  wire  _sum_T_1380 = sum_657 ^ sum_658; // @[Mul.scala 191:34]
  wire  sum_765 = sum_657 ^ sum_658 ^ cout_656; // @[Mul.scala 191:42]
  wire  cout_765 = sum_657 & sum_658 | _sum_T_1380 & cout_656; // @[Mul.scala 192:44]
  wire  sum_766 = sum_659 ^ sum_660; // @[Mul.scala 206:34]
  wire  cout_766 = sum_659 & sum_660; // @[Mul.scala 207:34]
  wire  sum_767 = cout_657 ^ cout_658; // @[Mul.scala 206:34]
  wire  cout_767 = cout_657 & cout_658; // @[Mul.scala 207:34]
  wire  sum_768 = sum_661 ^ sum_662; // @[Mul.scala 206:34]
  wire  cout_768 = sum_661 & sum_662; // @[Mul.scala 207:34]
  wire  sum_769 = cout_659 ^ cout_660; // @[Mul.scala 206:34]
  wire  cout_769 = cout_659 & cout_660; // @[Mul.scala 207:34]
  wire  sum_770 = sum_663 ^ sum_664; // @[Mul.scala 206:34]
  wire  cout_770 = sum_663 & sum_664; // @[Mul.scala 207:34]
  wire  sum_771 = cout_661 ^ cout_662; // @[Mul.scala 206:34]
  wire  cout_771 = cout_661 & cout_662; // @[Mul.scala 207:34]
  wire  sum_772 = sum_665 ^ sum_666; // @[Mul.scala 206:34]
  wire  cout_772 = sum_665 & sum_666; // @[Mul.scala 207:34]
  wire  sum_773 = cout_663 ^ cout_664; // @[Mul.scala 206:34]
  wire  cout_773 = cout_663 & cout_664; // @[Mul.scala 207:34]
  wire  sum_774 = sum_667 ^ sum_668; // @[Mul.scala 206:34]
  wire  cout_774 = sum_667 & sum_668; // @[Mul.scala 207:34]
  wire  sum_775 = cout_665 ^ cout_666; // @[Mul.scala 206:34]
  wire  cout_775 = cout_665 & cout_666; // @[Mul.scala 207:34]
  wire  sum_776 = sum_669 ^ sum_670; // @[Mul.scala 206:34]
  wire  cout_776 = sum_669 & sum_670; // @[Mul.scala 207:34]
  wire  sum_777 = cout_667 ^ cout_668; // @[Mul.scala 206:34]
  wire  cout_777 = cout_667 & cout_668; // @[Mul.scala 207:34]
  wire  sum_778 = sum_671 ^ sum_672; // @[Mul.scala 206:34]
  wire  cout_778 = sum_671 & sum_672; // @[Mul.scala 207:34]
  wire  sum_779 = cout_669 ^ cout_670; // @[Mul.scala 206:34]
  wire  cout_779 = cout_669 & cout_670; // @[Mul.scala 207:34]
  wire  sum_780 = sum_673 ^ sum_674; // @[Mul.scala 206:34]
  wire  cout_780 = sum_673 & sum_674; // @[Mul.scala 207:34]
  wire  sum_781 = cout_671 ^ cout_672; // @[Mul.scala 206:34]
  wire  cout_781 = cout_671 & cout_672; // @[Mul.scala 207:34]
  wire  sum_782 = sum_675 ^ sum_676; // @[Mul.scala 206:34]
  wire  cout_782 = sum_675 & sum_676; // @[Mul.scala 207:34]
  wire  sum_783 = cout_673 ^ cout_674; // @[Mul.scala 206:34]
  wire  cout_783 = cout_673 & cout_674; // @[Mul.scala 207:34]
  wire  sum_784 = sum_677 ^ sum_678; // @[Mul.scala 206:34]
  wire  cout_784 = sum_677 & sum_678; // @[Mul.scala 207:34]
  wire  sum_785 = cout_675 ^ cout_676; // @[Mul.scala 206:34]
  wire  cout_785 = cout_675 & cout_676; // @[Mul.scala 207:34]
  wire  sum_786 = sum_679 ^ sum_680; // @[Mul.scala 206:34]
  wire  cout_786 = sum_679 & sum_680; // @[Mul.scala 207:34]
  wire  sum_787 = cout_677 ^ cout_678; // @[Mul.scala 206:34]
  wire  cout_787 = cout_677 & cout_678; // @[Mul.scala 207:34]
  wire  sum_788 = sum_681 ^ sum_682; // @[Mul.scala 206:34]
  wire  cout_788 = sum_681 & sum_682; // @[Mul.scala 207:34]
  wire  sum_789 = cout_679 ^ cout_680; // @[Mul.scala 206:34]
  wire  cout_789 = cout_679 & cout_680; // @[Mul.scala 207:34]
  wire  sum_790 = sum_683 ^ sum_684; // @[Mul.scala 206:34]
  wire  cout_790 = sum_683 & sum_684; // @[Mul.scala 207:34]
  wire  sum_791 = cout_681 ^ cout_682; // @[Mul.scala 206:34]
  wire  cout_791 = cout_681 & cout_682; // @[Mul.scala 207:34]
  wire  sum_792 = sum_685 ^ sum_686; // @[Mul.scala 206:34]
  wire  cout_792 = sum_685 & sum_686; // @[Mul.scala 207:34]
  wire  sum_793 = cout_683 ^ cout_684; // @[Mul.scala 206:34]
  wire  cout_793 = cout_683 & cout_684; // @[Mul.scala 207:34]
  wire  sum_794 = sum_687 ^ sum_688; // @[Mul.scala 206:34]
  wire  cout_794 = sum_687 & sum_688; // @[Mul.scala 207:34]
  wire  sum_795 = cout_685 ^ cout_686; // @[Mul.scala 206:34]
  wire  cout_795 = cout_685 & cout_686; // @[Mul.scala 207:34]
  wire  sum_796 = sum_689 ^ sum_690; // @[Mul.scala 206:34]
  wire  cout_796 = sum_689 & sum_690; // @[Mul.scala 207:34]
  wire  sum_797 = cout_687 ^ cout_688; // @[Mul.scala 206:34]
  wire  cout_797 = cout_687 & cout_688; // @[Mul.scala 207:34]
  wire  sum_798 = sum_691 ^ sum_692; // @[Mul.scala 206:34]
  wire  cout_798 = sum_691 & sum_692; // @[Mul.scala 207:34]
  wire  sum_799 = cout_689 ^ cout_690; // @[Mul.scala 206:34]
  wire  cout_799 = cout_689 & cout_690; // @[Mul.scala 207:34]
  wire  sum_800 = sum_693 ^ sum_694; // @[Mul.scala 206:34]
  wire  cout_800 = sum_693 & sum_694; // @[Mul.scala 207:34]
  wire  sum_801 = cout_691 ^ cout_692; // @[Mul.scala 206:34]
  wire  cout_801 = cout_691 & cout_692; // @[Mul.scala 207:34]
  wire  sum_802 = sum_695 ^ sum_696; // @[Mul.scala 206:34]
  wire  cout_802 = sum_695 & sum_696; // @[Mul.scala 207:34]
  wire  sum_803 = cout_693 ^ cout_694; // @[Mul.scala 206:34]
  wire  cout_803 = cout_693 & cout_694; // @[Mul.scala 207:34]
  wire  sum_804 = sum_697 ^ sum_698; // @[Mul.scala 206:34]
  wire  cout_804 = sum_697 & sum_698; // @[Mul.scala 207:34]
  wire  sum_805 = cout_695 ^ cout_696; // @[Mul.scala 206:34]
  wire  cout_805 = cout_695 & cout_696; // @[Mul.scala 207:34]
  wire  sum_806 = sum_699 ^ sum_700; // @[Mul.scala 206:34]
  wire  cout_806 = sum_699 & sum_700; // @[Mul.scala 207:34]
  wire  sum_807 = cout_697 ^ cout_698; // @[Mul.scala 206:34]
  wire  cout_807 = cout_697 & cout_698; // @[Mul.scala 207:34]
  wire  sum_808 = sum_701 ^ sum_702; // @[Mul.scala 206:34]
  wire  cout_808 = sum_701 & sum_702; // @[Mul.scala 207:34]
  wire  sum_809 = cout_699 ^ cout_700; // @[Mul.scala 206:34]
  wire  cout_809 = cout_699 & cout_700; // @[Mul.scala 207:34]
  wire  sum_810 = sum_703 ^ sum_704; // @[Mul.scala 206:34]
  wire  cout_810 = sum_703 & sum_704; // @[Mul.scala 207:34]
  wire  sum_811 = cout_701 ^ cout_702; // @[Mul.scala 206:34]
  wire  cout_811 = cout_701 & cout_702; // @[Mul.scala 207:34]
  wire  sum_812 = sum_705 ^ sum_706; // @[Mul.scala 206:34]
  wire  cout_812 = sum_705 & sum_706; // @[Mul.scala 207:34]
  wire  sum_813 = cout_703 ^ cout_704; // @[Mul.scala 206:34]
  wire  cout_813 = cout_703 & cout_704; // @[Mul.scala 207:34]
  wire  sum_814 = sum_707 ^ sum_708; // @[Mul.scala 206:34]
  wire  cout_814 = sum_707 & sum_708; // @[Mul.scala 207:34]
  wire  sum_815 = cout_705 ^ cout_706; // @[Mul.scala 206:34]
  wire  cout_815 = cout_705 & cout_706; // @[Mul.scala 207:34]
  wire  sum_816 = sum_709 ^ sum_710; // @[Mul.scala 206:34]
  wire  cout_816 = sum_709 & sum_710; // @[Mul.scala 207:34]
  wire  sum_817 = cout_707 ^ cout_708; // @[Mul.scala 206:34]
  wire  cout_817 = cout_707 & cout_708; // @[Mul.scala 207:34]
  wire  sum_818 = sum_711 ^ sum_712; // @[Mul.scala 206:34]
  wire  cout_818 = sum_711 & sum_712; // @[Mul.scala 207:34]
  wire  sum_819 = cout_709 ^ cout_710; // @[Mul.scala 206:34]
  wire  cout_819 = cout_709 & cout_710; // @[Mul.scala 207:34]
  wire  sum_820 = sum_713 ^ sum_714; // @[Mul.scala 206:34]
  wire  cout_820 = sum_713 & sum_714; // @[Mul.scala 207:34]
  wire  sum_821 = cout_711 ^ cout_712; // @[Mul.scala 206:34]
  wire  cout_821 = cout_711 & cout_712; // @[Mul.scala 207:34]
  wire  sum_822 = sum_715 ^ sum_716; // @[Mul.scala 206:34]
  wire  cout_822 = sum_715 & sum_716; // @[Mul.scala 207:34]
  wire  sum_823 = cout_713 ^ cout_714; // @[Mul.scala 206:34]
  wire  cout_823 = cout_713 & cout_714; // @[Mul.scala 207:34]
  wire  sum_824 = sum_717 ^ sum_718; // @[Mul.scala 206:34]
  wire  cout_824 = sum_717 & sum_718; // @[Mul.scala 207:34]
  wire  sum_825 = cout_715 ^ cout_716; // @[Mul.scala 206:34]
  wire  cout_825 = cout_715 & cout_716; // @[Mul.scala 207:34]
  wire  sum_826 = sum_719 ^ sum_720; // @[Mul.scala 206:34]
  wire  cout_826 = sum_719 & sum_720; // @[Mul.scala 207:34]
  wire  sum_827 = cout_717 ^ cout_718; // @[Mul.scala 206:34]
  wire  cout_827 = cout_717 & cout_718; // @[Mul.scala 207:34]
  wire  sum_828 = sum_721 ^ sum_722; // @[Mul.scala 206:34]
  wire  cout_828 = sum_721 & sum_722; // @[Mul.scala 207:34]
  wire  sum_829 = cout_719 ^ cout_720; // @[Mul.scala 206:34]
  wire  cout_829 = cout_719 & cout_720; // @[Mul.scala 207:34]
  wire  sum_830 = sum_723 ^ sum_724; // @[Mul.scala 206:34]
  wire  cout_830 = sum_723 & sum_724; // @[Mul.scala 207:34]
  wire  sum_831 = cout_721 ^ cout_722; // @[Mul.scala 206:34]
  wire  cout_831 = cout_721 & cout_722; // @[Mul.scala 207:34]
  wire  sum_832 = sum_725 ^ sum_726; // @[Mul.scala 206:34]
  wire  cout_832 = sum_725 & sum_726; // @[Mul.scala 207:34]
  wire  sum_833 = cout_723 ^ cout_724; // @[Mul.scala 206:34]
  wire  cout_833 = cout_723 & cout_724; // @[Mul.scala 207:34]
  wire  sum_834 = sum_727 ^ sum_728; // @[Mul.scala 206:34]
  wire  cout_834 = sum_727 & sum_728; // @[Mul.scala 207:34]
  wire  sum_835 = cout_725 ^ cout_726; // @[Mul.scala 206:34]
  wire  cout_835 = cout_725 & cout_726; // @[Mul.scala 207:34]
  wire  sum_836 = sum_729 ^ sum_730; // @[Mul.scala 206:34]
  wire  cout_836 = sum_729 & sum_730; // @[Mul.scala 207:34]
  wire  sum_837 = cout_727 ^ cout_728; // @[Mul.scala 206:34]
  wire  cout_837 = cout_727 & cout_728; // @[Mul.scala 207:34]
  wire  sum_838 = sum_731 ^ sum_732; // @[Mul.scala 206:34]
  wire  cout_838 = sum_731 & sum_732; // @[Mul.scala 207:34]
  wire  sum_839 = cout_729 ^ cout_730; // @[Mul.scala 206:34]
  wire  cout_839 = cout_729 & cout_730; // @[Mul.scala 207:34]
  wire  sum_840 = sum_733 ^ sum_734; // @[Mul.scala 206:34]
  wire  cout_840 = sum_733 & sum_734; // @[Mul.scala 207:34]
  wire  sum_841 = cout_731 ^ cout_732; // @[Mul.scala 206:34]
  wire  cout_841 = cout_731 & cout_732; // @[Mul.scala 207:34]
  wire  sum_842 = sum_735 ^ sum_736; // @[Mul.scala 206:34]
  wire  cout_842 = sum_735 & sum_736; // @[Mul.scala 207:34]
  wire  sum_843 = cout_733 ^ cout_734; // @[Mul.scala 206:34]
  wire  cout_843 = cout_733 & cout_734; // @[Mul.scala 207:34]
  wire  sum_844 = sum_737 ^ sum_738; // @[Mul.scala 206:34]
  wire  cout_844 = sum_737 & sum_738; // @[Mul.scala 207:34]
  wire  sum_845 = cout_735 ^ cout_736; // @[Mul.scala 206:34]
  wire  cout_845 = cout_735 & cout_736; // @[Mul.scala 207:34]
  wire  sum_846 = sum_739 ^ sum_740; // @[Mul.scala 206:34]
  wire  cout_846 = sum_739 & sum_740; // @[Mul.scala 207:34]
  wire  sum_847 = cout_737 ^ cout_738; // @[Mul.scala 206:34]
  wire  cout_847 = cout_737 & cout_738; // @[Mul.scala 207:34]
  wire  sum_848 = sum_741 ^ sum_742; // @[Mul.scala 206:34]
  wire  cout_848 = sum_741 & sum_742; // @[Mul.scala 207:34]
  wire  sum_849 = cout_739 ^ cout_740; // @[Mul.scala 206:34]
  wire  cout_849 = cout_739 & cout_740; // @[Mul.scala 207:34]
  wire  sum_850 = sum_743 ^ sum_744; // @[Mul.scala 206:34]
  wire  cout_850 = sum_743 & sum_744; // @[Mul.scala 207:34]
  wire  sum_851 = cout_741 ^ cout_742; // @[Mul.scala 206:34]
  wire  cout_851 = cout_741 & cout_742; // @[Mul.scala 207:34]
  wire  sum_852 = sum_745 ^ sum_746; // @[Mul.scala 206:34]
  wire  cout_852 = sum_745 & sum_746; // @[Mul.scala 207:34]
  wire  sum_853 = cout_743 ^ cout_744; // @[Mul.scala 206:34]
  wire  cout_853 = cout_743 & cout_744; // @[Mul.scala 207:34]
  wire  _sum_T_1470 = sum_747 ^ cout_745; // @[Mul.scala 191:34]
  wire  sum_854 = sum_747 ^ cout_745 ^ cout_746; // @[Mul.scala 191:42]
  wire  cout_854 = sum_747 & cout_745 | _sum_T_1470 & cout_746; // @[Mul.scala 192:44]
  wire  sum_855 = sum_748 ^ cout_747; // @[Mul.scala 206:34]
  wire  cout_855 = sum_748 & cout_747; // @[Mul.scala 207:34]
  wire  sum_856 = sum_749 ^ cout_748; // @[Mul.scala 206:34]
  wire  cout_856 = sum_749 & cout_748; // @[Mul.scala 207:34]
  wire  sum_857 = sum_750 ^ cout_749; // @[Mul.scala 206:34]
  wire  cout_857 = sum_750 & cout_749; // @[Mul.scala 207:34]
  wire  sum_858 = sum_751 ^ cout_750; // @[Mul.scala 206:34]
  wire  cout_858 = sum_751 & cout_750; // @[Mul.scala 207:34]
  wire  sum_859 = sum_752 ^ cout_751; // @[Mul.scala 206:34]
  wire  sum_870 = sum_763 ^ cout_762; // @[Mul.scala 206:34]
  wire  cout_870 = sum_763 & cout_762; // @[Mul.scala 207:34]
  wire  sum_871 = sum_764 ^ cout_763; // @[Mul.scala 206:34]
  wire  cout_871 = sum_764 & cout_763; // @[Mul.scala 207:34]
  wire  sum_872 = sum_765 ^ cout_764; // @[Mul.scala 206:34]
  wire  cout_872 = sum_765 & cout_764; // @[Mul.scala 207:34]
  wire  _sum_T_1490 = sum_766 ^ sum_767; // @[Mul.scala 191:34]
  wire  sum_873 = sum_766 ^ sum_767 ^ cout_765; // @[Mul.scala 191:42]
  wire  cout_873 = sum_766 & sum_767 | _sum_T_1490 & cout_765; // @[Mul.scala 192:44]
  wire  sum_874 = sum_768 ^ sum_769; // @[Mul.scala 206:34]
  wire  cout_874 = sum_768 & sum_769; // @[Mul.scala 207:34]
  wire  sum_875 = cout_766 ^ cout_767; // @[Mul.scala 206:34]
  wire  cout_875 = cout_766 & cout_767; // @[Mul.scala 207:34]
  wire  sum_876 = sum_770 ^ sum_771; // @[Mul.scala 206:34]
  wire  cout_876 = sum_770 & sum_771; // @[Mul.scala 207:34]
  wire  sum_877 = cout_768 ^ cout_769; // @[Mul.scala 206:34]
  wire  cout_877 = cout_768 & cout_769; // @[Mul.scala 207:34]
  wire  sum_878 = sum_772 ^ sum_773; // @[Mul.scala 206:34]
  wire  cout_878 = sum_772 & sum_773; // @[Mul.scala 207:34]
  wire  sum_879 = cout_770 ^ cout_771; // @[Mul.scala 206:34]
  wire  cout_879 = cout_770 & cout_771; // @[Mul.scala 207:34]
  wire  sum_880 = sum_774 ^ sum_775; // @[Mul.scala 206:34]
  wire  cout_880 = sum_774 & sum_775; // @[Mul.scala 207:34]
  wire  sum_881 = cout_772 ^ cout_773; // @[Mul.scala 206:34]
  wire  cout_881 = cout_772 & cout_773; // @[Mul.scala 207:34]
  wire  sum_882 = sum_776 ^ sum_777; // @[Mul.scala 206:34]
  wire  cout_882 = sum_776 & sum_777; // @[Mul.scala 207:34]
  wire  sum_883 = cout_774 ^ cout_775; // @[Mul.scala 206:34]
  wire  cout_883 = cout_774 & cout_775; // @[Mul.scala 207:34]
  wire  sum_884 = sum_778 ^ sum_779; // @[Mul.scala 206:34]
  wire  cout_884 = sum_778 & sum_779; // @[Mul.scala 207:34]
  wire  sum_885 = cout_776 ^ cout_777; // @[Mul.scala 206:34]
  wire  cout_885 = cout_776 & cout_777; // @[Mul.scala 207:34]
  wire  sum_886 = sum_780 ^ sum_781; // @[Mul.scala 206:34]
  wire  cout_886 = sum_780 & sum_781; // @[Mul.scala 207:34]
  wire  sum_887 = cout_778 ^ cout_779; // @[Mul.scala 206:34]
  wire  cout_887 = cout_778 & cout_779; // @[Mul.scala 207:34]
  wire  sum_888 = sum_782 ^ sum_783; // @[Mul.scala 206:34]
  wire  cout_888 = sum_782 & sum_783; // @[Mul.scala 207:34]
  wire  sum_889 = cout_780 ^ cout_781; // @[Mul.scala 206:34]
  wire  cout_889 = cout_780 & cout_781; // @[Mul.scala 207:34]
  wire  sum_890 = sum_784 ^ sum_785; // @[Mul.scala 206:34]
  wire  cout_890 = sum_784 & sum_785; // @[Mul.scala 207:34]
  wire  sum_891 = cout_782 ^ cout_783; // @[Mul.scala 206:34]
  wire  cout_891 = cout_782 & cout_783; // @[Mul.scala 207:34]
  wire  sum_892 = sum_786 ^ sum_787; // @[Mul.scala 206:34]
  wire  cout_892 = sum_786 & sum_787; // @[Mul.scala 207:34]
  wire  sum_893 = cout_784 ^ cout_785; // @[Mul.scala 206:34]
  wire  cout_893 = cout_784 & cout_785; // @[Mul.scala 207:34]
  wire  sum_894 = sum_788 ^ sum_789; // @[Mul.scala 206:34]
  wire  cout_894 = sum_788 & sum_789; // @[Mul.scala 207:34]
  wire  sum_895 = cout_786 ^ cout_787; // @[Mul.scala 206:34]
  wire  cout_895 = cout_786 & cout_787; // @[Mul.scala 207:34]
  wire  sum_896 = sum_790 ^ sum_791; // @[Mul.scala 206:34]
  wire  cout_896 = sum_790 & sum_791; // @[Mul.scala 207:34]
  wire  sum_897 = cout_788 ^ cout_789; // @[Mul.scala 206:34]
  wire  cout_897 = cout_788 & cout_789; // @[Mul.scala 207:34]
  wire  sum_898 = sum_792 ^ sum_793; // @[Mul.scala 206:34]
  wire  cout_898 = sum_792 & sum_793; // @[Mul.scala 207:34]
  wire  sum_899 = cout_790 ^ cout_791; // @[Mul.scala 206:34]
  wire  cout_899 = cout_790 & cout_791; // @[Mul.scala 207:34]
  wire  sum_900 = sum_794 ^ sum_795; // @[Mul.scala 206:34]
  wire  cout_900 = sum_794 & sum_795; // @[Mul.scala 207:34]
  wire  sum_901 = cout_792 ^ cout_793; // @[Mul.scala 206:34]
  wire  cout_901 = cout_792 & cout_793; // @[Mul.scala 207:34]
  wire  sum_902 = sum_796 ^ sum_797; // @[Mul.scala 206:34]
  wire  cout_902 = sum_796 & sum_797; // @[Mul.scala 207:34]
  wire  sum_903 = cout_794 ^ cout_795; // @[Mul.scala 206:34]
  wire  cout_903 = cout_794 & cout_795; // @[Mul.scala 207:34]
  wire  sum_904 = sum_798 ^ sum_799; // @[Mul.scala 206:34]
  wire  cout_904 = sum_798 & sum_799; // @[Mul.scala 207:34]
  wire  sum_905 = cout_796 ^ cout_797; // @[Mul.scala 206:34]
  wire  cout_905 = cout_796 & cout_797; // @[Mul.scala 207:34]
  wire  sum_906 = sum_800 ^ sum_801; // @[Mul.scala 206:34]
  wire  cout_906 = sum_800 & sum_801; // @[Mul.scala 207:34]
  wire  sum_907 = cout_798 ^ cout_799; // @[Mul.scala 206:34]
  wire  cout_907 = cout_798 & cout_799; // @[Mul.scala 207:34]
  wire  sum_908 = sum_802 ^ sum_803; // @[Mul.scala 206:34]
  wire  cout_908 = sum_802 & sum_803; // @[Mul.scala 207:34]
  wire  sum_909 = cout_800 ^ cout_801; // @[Mul.scala 206:34]
  wire  cout_909 = cout_800 & cout_801; // @[Mul.scala 207:34]
  wire  sum_910 = sum_804 ^ sum_805; // @[Mul.scala 206:34]
  wire  cout_910 = sum_804 & sum_805; // @[Mul.scala 207:34]
  wire  sum_911 = cout_802 ^ cout_803; // @[Mul.scala 206:34]
  wire  cout_911 = cout_802 & cout_803; // @[Mul.scala 207:34]
  wire  sum_912 = sum_806 ^ sum_807; // @[Mul.scala 206:34]
  wire  cout_912 = sum_806 & sum_807; // @[Mul.scala 207:34]
  wire  sum_913 = cout_804 ^ cout_805; // @[Mul.scala 206:34]
  wire  cout_913 = cout_804 & cout_805; // @[Mul.scala 207:34]
  wire  sum_914 = sum_808 ^ sum_809; // @[Mul.scala 206:34]
  wire  cout_914 = sum_808 & sum_809; // @[Mul.scala 207:34]
  wire  sum_915 = cout_806 ^ cout_807; // @[Mul.scala 206:34]
  wire  cout_915 = cout_806 & cout_807; // @[Mul.scala 207:34]
  wire  sum_916 = sum_810 ^ sum_811; // @[Mul.scala 206:34]
  wire  cout_916 = sum_810 & sum_811; // @[Mul.scala 207:34]
  wire  sum_917 = cout_808 ^ cout_809; // @[Mul.scala 206:34]
  wire  cout_917 = cout_808 & cout_809; // @[Mul.scala 207:34]
  wire  sum_918 = sum_812 ^ sum_813; // @[Mul.scala 206:34]
  wire  cout_918 = sum_812 & sum_813; // @[Mul.scala 207:34]
  wire  sum_919 = cout_810 ^ cout_811; // @[Mul.scala 206:34]
  wire  cout_919 = cout_810 & cout_811; // @[Mul.scala 207:34]
  wire  sum_920 = sum_814 ^ sum_815; // @[Mul.scala 206:34]
  wire  cout_920 = sum_814 & sum_815; // @[Mul.scala 207:34]
  wire  sum_921 = cout_812 ^ cout_813; // @[Mul.scala 206:34]
  wire  cout_921 = cout_812 & cout_813; // @[Mul.scala 207:34]
  wire  sum_922 = sum_816 ^ sum_817; // @[Mul.scala 206:34]
  wire  cout_922 = sum_816 & sum_817; // @[Mul.scala 207:34]
  wire  sum_923 = cout_814 ^ cout_815; // @[Mul.scala 206:34]
  wire  cout_923 = cout_814 & cout_815; // @[Mul.scala 207:34]
  wire  sum_924 = sum_818 ^ sum_819; // @[Mul.scala 206:34]
  wire  cout_924 = sum_818 & sum_819; // @[Mul.scala 207:34]
  wire  sum_925 = cout_816 ^ cout_817; // @[Mul.scala 206:34]
  wire  cout_925 = cout_816 & cout_817; // @[Mul.scala 207:34]
  wire  sum_926 = sum_820 ^ sum_821; // @[Mul.scala 206:34]
  wire  cout_926 = sum_820 & sum_821; // @[Mul.scala 207:34]
  wire  sum_927 = cout_818 ^ cout_819; // @[Mul.scala 206:34]
  wire  cout_927 = cout_818 & cout_819; // @[Mul.scala 207:34]
  wire  sum_928 = sum_822 ^ sum_823; // @[Mul.scala 206:34]
  wire  cout_928 = sum_822 & sum_823; // @[Mul.scala 207:34]
  wire  sum_929 = cout_820 ^ cout_821; // @[Mul.scala 206:34]
  wire  cout_929 = cout_820 & cout_821; // @[Mul.scala 207:34]
  wire  sum_930 = sum_824 ^ sum_825; // @[Mul.scala 206:34]
  wire  cout_930 = sum_824 & sum_825; // @[Mul.scala 207:34]
  wire  sum_931 = cout_822 ^ cout_823; // @[Mul.scala 206:34]
  wire  cout_931 = cout_822 & cout_823; // @[Mul.scala 207:34]
  wire  sum_932 = sum_826 ^ sum_827; // @[Mul.scala 206:34]
  wire  cout_932 = sum_826 & sum_827; // @[Mul.scala 207:34]
  wire  sum_933 = cout_824 ^ cout_825; // @[Mul.scala 206:34]
  wire  cout_933 = cout_824 & cout_825; // @[Mul.scala 207:34]
  wire  sum_934 = sum_828 ^ sum_829; // @[Mul.scala 206:34]
  wire  cout_934 = sum_828 & sum_829; // @[Mul.scala 207:34]
  wire  sum_935 = cout_826 ^ cout_827; // @[Mul.scala 206:34]
  wire  cout_935 = cout_826 & cout_827; // @[Mul.scala 207:34]
  wire  sum_936 = sum_830 ^ sum_831; // @[Mul.scala 206:34]
  wire  cout_936 = sum_830 & sum_831; // @[Mul.scala 207:34]
  wire  sum_937 = cout_828 ^ cout_829; // @[Mul.scala 206:34]
  wire  cout_937 = cout_828 & cout_829; // @[Mul.scala 207:34]
  wire  sum_938 = sum_832 ^ sum_833; // @[Mul.scala 206:34]
  wire  cout_938 = sum_832 & sum_833; // @[Mul.scala 207:34]
  wire  sum_939 = cout_830 ^ cout_831; // @[Mul.scala 206:34]
  wire  cout_939 = cout_830 & cout_831; // @[Mul.scala 207:34]
  wire  sum_940 = sum_834 ^ sum_835; // @[Mul.scala 206:34]
  wire  cout_940 = sum_834 & sum_835; // @[Mul.scala 207:34]
  wire  sum_941 = cout_832 ^ cout_833; // @[Mul.scala 206:34]
  wire  cout_941 = cout_832 & cout_833; // @[Mul.scala 207:34]
  wire  sum_942 = sum_836 ^ sum_837; // @[Mul.scala 206:34]
  wire  cout_942 = sum_836 & sum_837; // @[Mul.scala 207:34]
  wire  sum_943 = cout_834 ^ cout_835; // @[Mul.scala 206:34]
  wire  cout_943 = cout_834 & cout_835; // @[Mul.scala 207:34]
  wire  sum_944 = sum_838 ^ sum_839; // @[Mul.scala 206:34]
  wire  cout_944 = sum_838 & sum_839; // @[Mul.scala 207:34]
  wire  sum_945 = cout_836 ^ cout_837; // @[Mul.scala 206:34]
  wire  cout_945 = cout_836 & cout_837; // @[Mul.scala 207:34]
  wire  sum_946 = sum_840 ^ sum_841; // @[Mul.scala 206:34]
  wire  cout_946 = sum_840 & sum_841; // @[Mul.scala 207:34]
  wire  sum_947 = cout_838 ^ cout_839; // @[Mul.scala 206:34]
  wire  cout_947 = cout_838 & cout_839; // @[Mul.scala 207:34]
  wire  sum_948 = sum_842 ^ sum_843; // @[Mul.scala 206:34]
  wire  cout_948 = sum_842 & sum_843; // @[Mul.scala 207:34]
  wire  sum_949 = cout_840 ^ cout_841; // @[Mul.scala 206:34]
  wire  cout_949 = cout_840 & cout_841; // @[Mul.scala 207:34]
  wire  sum_950 = sum_844 ^ sum_845; // @[Mul.scala 206:34]
  wire  cout_950 = sum_844 & sum_845; // @[Mul.scala 207:34]
  wire  sum_951 = cout_842 ^ cout_843; // @[Mul.scala 206:34]
  wire  cout_951 = cout_842 & cout_843; // @[Mul.scala 207:34]
  wire  sum_952 = sum_846 ^ sum_847; // @[Mul.scala 206:34]
  wire  cout_952 = sum_846 & sum_847; // @[Mul.scala 207:34]
  wire  sum_953 = cout_844 ^ cout_845; // @[Mul.scala 206:34]
  wire  cout_953 = cout_844 & cout_845; // @[Mul.scala 207:34]
  wire  sum_954 = sum_848 ^ sum_849; // @[Mul.scala 206:34]
  wire  cout_954 = sum_848 & sum_849; // @[Mul.scala 207:34]
  wire  sum_955 = cout_846 ^ cout_847; // @[Mul.scala 206:34]
  wire  cout_955 = cout_846 & cout_847; // @[Mul.scala 207:34]
  wire  sum_956 = sum_850 ^ sum_851; // @[Mul.scala 206:34]
  wire  cout_956 = sum_850 & sum_851; // @[Mul.scala 207:34]
  wire  sum_957 = cout_848 ^ cout_849; // @[Mul.scala 206:34]
  wire  cout_957 = cout_848 & cout_849; // @[Mul.scala 207:34]
  wire  sum_958 = sum_852 ^ sum_853; // @[Mul.scala 206:34]
  wire  cout_958 = sum_852 & sum_853; // @[Mul.scala 207:34]
  wire  sum_959 = cout_850 ^ cout_851; // @[Mul.scala 206:34]
  wire  cout_959 = cout_850 & cout_851; // @[Mul.scala 207:34]
  wire  _sum_T_1578 = sum_854 ^ cout_852; // @[Mul.scala 191:34]
  wire  sum_960 = sum_854 ^ cout_852 ^ cout_853; // @[Mul.scala 191:42]
  wire  cout_960 = sum_854 & cout_852 | _sum_T_1578 & cout_853; // @[Mul.scala 192:44]
  wire  sum_961 = sum_855 ^ cout_854; // @[Mul.scala 206:34]
  wire  cout_961 = sum_855 & cout_854; // @[Mul.scala 207:34]
  wire  sum_962 = sum_856 ^ cout_855; // @[Mul.scala 206:34]
  wire  cout_962 = sum_856 & cout_855; // @[Mul.scala 207:34]
  wire  sum_963 = sum_857 ^ cout_856; // @[Mul.scala 206:34]
  wire  cout_963 = sum_857 & cout_856; // @[Mul.scala 207:34]
  wire  sum_964 = sum_858 ^ cout_857; // @[Mul.scala 206:34]
  wire  cout_964 = sum_858 & cout_857; // @[Mul.scala 207:34]
  wire  sum_965 = sum_859 ^ cout_858; // @[Mul.scala 206:34]
  wire  sum_977 = sum_871 ^ cout_870; // @[Mul.scala 206:34]
  wire  cout_977 = sum_871 & cout_870; // @[Mul.scala 207:34]
  wire  sum_978 = sum_872 ^ cout_871; // @[Mul.scala 206:34]
  wire  cout_978 = sum_872 & cout_871; // @[Mul.scala 207:34]
  wire  sum_979 = sum_873 ^ cout_872; // @[Mul.scala 206:34]
  wire  cout_979 = sum_873 & cout_872; // @[Mul.scala 207:34]
  wire  _sum_T_1599 = sum_874 ^ sum_875; // @[Mul.scala 191:34]
  wire  sum_980 = sum_874 ^ sum_875 ^ cout_873; // @[Mul.scala 191:42]
  wire  cout_980 = sum_874 & sum_875 | _sum_T_1599 & cout_873; // @[Mul.scala 192:44]
  wire  sum_981 = sum_876 ^ sum_877; // @[Mul.scala 206:34]
  wire  cout_981 = sum_876 & sum_877; // @[Mul.scala 207:34]
  wire  sum_982 = cout_874 ^ cout_875; // @[Mul.scala 206:34]
  wire  cout_982 = cout_874 & cout_875; // @[Mul.scala 207:34]
  wire  sum_983 = sum_878 ^ sum_879; // @[Mul.scala 206:34]
  wire  cout_983 = sum_878 & sum_879; // @[Mul.scala 207:34]
  wire  sum_984 = cout_876 ^ cout_877; // @[Mul.scala 206:34]
  wire  cout_984 = cout_876 & cout_877; // @[Mul.scala 207:34]
  wire  sum_985 = sum_880 ^ sum_881; // @[Mul.scala 206:34]
  wire  cout_985 = sum_880 & sum_881; // @[Mul.scala 207:34]
  wire  sum_986 = cout_878 ^ cout_879; // @[Mul.scala 206:34]
  wire  cout_986 = cout_878 & cout_879; // @[Mul.scala 207:34]
  wire  sum_987 = sum_882 ^ sum_883; // @[Mul.scala 206:34]
  wire  cout_987 = sum_882 & sum_883; // @[Mul.scala 207:34]
  wire  sum_988 = cout_880 ^ cout_881; // @[Mul.scala 206:34]
  wire  cout_988 = cout_880 & cout_881; // @[Mul.scala 207:34]
  wire  sum_989 = sum_884 ^ sum_885; // @[Mul.scala 206:34]
  wire  cout_989 = sum_884 & sum_885; // @[Mul.scala 207:34]
  wire  sum_990 = cout_882 ^ cout_883; // @[Mul.scala 206:34]
  wire  cout_990 = cout_882 & cout_883; // @[Mul.scala 207:34]
  wire  sum_991 = sum_886 ^ sum_887; // @[Mul.scala 206:34]
  wire  cout_991 = sum_886 & sum_887; // @[Mul.scala 207:34]
  wire  sum_992 = cout_884 ^ cout_885; // @[Mul.scala 206:34]
  wire  cout_992 = cout_884 & cout_885; // @[Mul.scala 207:34]
  wire  sum_993 = sum_888 ^ sum_889; // @[Mul.scala 206:34]
  wire  cout_993 = sum_888 & sum_889; // @[Mul.scala 207:34]
  wire  sum_994 = cout_886 ^ cout_887; // @[Mul.scala 206:34]
  wire  cout_994 = cout_886 & cout_887; // @[Mul.scala 207:34]
  wire  sum_995 = sum_890 ^ sum_891; // @[Mul.scala 206:34]
  wire  cout_995 = sum_890 & sum_891; // @[Mul.scala 207:34]
  wire  sum_996 = cout_888 ^ cout_889; // @[Mul.scala 206:34]
  wire  cout_996 = cout_888 & cout_889; // @[Mul.scala 207:34]
  wire  sum_997 = sum_892 ^ sum_893; // @[Mul.scala 206:34]
  wire  cout_997 = sum_892 & sum_893; // @[Mul.scala 207:34]
  wire  sum_998 = cout_890 ^ cout_891; // @[Mul.scala 206:34]
  wire  cout_998 = cout_890 & cout_891; // @[Mul.scala 207:34]
  wire  sum_999 = sum_894 ^ sum_895; // @[Mul.scala 206:34]
  wire  cout_999 = sum_894 & sum_895; // @[Mul.scala 207:34]
  wire  sum_1000 = cout_892 ^ cout_893; // @[Mul.scala 206:34]
  wire  cout_1000 = cout_892 & cout_893; // @[Mul.scala 207:34]
  wire  sum_1001 = sum_896 ^ sum_897; // @[Mul.scala 206:34]
  wire  cout_1001 = sum_896 & sum_897; // @[Mul.scala 207:34]
  wire  sum_1002 = cout_894 ^ cout_895; // @[Mul.scala 206:34]
  wire  cout_1002 = cout_894 & cout_895; // @[Mul.scala 207:34]
  wire  sum_1003 = sum_898 ^ sum_899; // @[Mul.scala 206:34]
  wire  cout_1003 = sum_898 & sum_899; // @[Mul.scala 207:34]
  wire  sum_1004 = cout_896 ^ cout_897; // @[Mul.scala 206:34]
  wire  cout_1004 = cout_896 & cout_897; // @[Mul.scala 207:34]
  wire  sum_1005 = sum_900 ^ sum_901; // @[Mul.scala 206:34]
  wire  cout_1005 = sum_900 & sum_901; // @[Mul.scala 207:34]
  wire  sum_1006 = cout_898 ^ cout_899; // @[Mul.scala 206:34]
  wire  cout_1006 = cout_898 & cout_899; // @[Mul.scala 207:34]
  wire  sum_1007 = sum_902 ^ sum_903; // @[Mul.scala 206:34]
  wire  cout_1007 = sum_902 & sum_903; // @[Mul.scala 207:34]
  wire  sum_1008 = cout_900 ^ cout_901; // @[Mul.scala 206:34]
  wire  cout_1008 = cout_900 & cout_901; // @[Mul.scala 207:34]
  wire  sum_1009 = sum_904 ^ sum_905; // @[Mul.scala 206:34]
  wire  cout_1009 = sum_904 & sum_905; // @[Mul.scala 207:34]
  wire  sum_1010 = cout_902 ^ cout_903; // @[Mul.scala 206:34]
  wire  cout_1010 = cout_902 & cout_903; // @[Mul.scala 207:34]
  wire  sum_1011 = sum_906 ^ sum_907; // @[Mul.scala 206:34]
  wire  cout_1011 = sum_906 & sum_907; // @[Mul.scala 207:34]
  wire  sum_1012 = cout_904 ^ cout_905; // @[Mul.scala 206:34]
  wire  cout_1012 = cout_904 & cout_905; // @[Mul.scala 207:34]
  wire  sum_1013 = sum_908 ^ sum_909; // @[Mul.scala 206:34]
  wire  cout_1013 = sum_908 & sum_909; // @[Mul.scala 207:34]
  wire  sum_1014 = cout_906 ^ cout_907; // @[Mul.scala 206:34]
  wire  cout_1014 = cout_906 & cout_907; // @[Mul.scala 207:34]
  wire  sum_1015 = sum_910 ^ sum_911; // @[Mul.scala 206:34]
  wire  cout_1015 = sum_910 & sum_911; // @[Mul.scala 207:34]
  wire  sum_1016 = cout_908 ^ cout_909; // @[Mul.scala 206:34]
  wire  cout_1016 = cout_908 & cout_909; // @[Mul.scala 207:34]
  wire  sum_1017 = sum_912 ^ sum_913; // @[Mul.scala 206:34]
  wire  cout_1017 = sum_912 & sum_913; // @[Mul.scala 207:34]
  wire  sum_1018 = cout_910 ^ cout_911; // @[Mul.scala 206:34]
  wire  cout_1018 = cout_910 & cout_911; // @[Mul.scala 207:34]
  wire  sum_1019 = sum_914 ^ sum_915; // @[Mul.scala 206:34]
  wire  cout_1019 = sum_914 & sum_915; // @[Mul.scala 207:34]
  wire  sum_1020 = cout_912 ^ cout_913; // @[Mul.scala 206:34]
  wire  cout_1020 = cout_912 & cout_913; // @[Mul.scala 207:34]
  wire  sum_1021 = sum_916 ^ sum_917; // @[Mul.scala 206:34]
  wire  cout_1021 = sum_916 & sum_917; // @[Mul.scala 207:34]
  wire  sum_1022 = cout_914 ^ cout_915; // @[Mul.scala 206:34]
  wire  cout_1022 = cout_914 & cout_915; // @[Mul.scala 207:34]
  wire  sum_1023 = sum_918 ^ sum_919; // @[Mul.scala 206:34]
  wire  cout_1023 = sum_918 & sum_919; // @[Mul.scala 207:34]
  wire  sum_1024 = cout_916 ^ cout_917; // @[Mul.scala 206:34]
  wire  cout_1024 = cout_916 & cout_917; // @[Mul.scala 207:34]
  wire  sum_1025 = sum_920 ^ sum_921; // @[Mul.scala 206:34]
  wire  cout_1025 = sum_920 & sum_921; // @[Mul.scala 207:34]
  wire  sum_1026 = cout_918 ^ cout_919; // @[Mul.scala 206:34]
  wire  cout_1026 = cout_918 & cout_919; // @[Mul.scala 207:34]
  wire  sum_1027 = sum_922 ^ sum_923; // @[Mul.scala 206:34]
  wire  cout_1027 = sum_922 & sum_923; // @[Mul.scala 207:34]
  wire  sum_1028 = cout_920 ^ cout_921; // @[Mul.scala 206:34]
  wire  cout_1028 = cout_920 & cout_921; // @[Mul.scala 207:34]
  wire  sum_1029 = sum_924 ^ sum_925; // @[Mul.scala 206:34]
  wire  cout_1029 = sum_924 & sum_925; // @[Mul.scala 207:34]
  wire  sum_1030 = cout_922 ^ cout_923; // @[Mul.scala 206:34]
  wire  cout_1030 = cout_922 & cout_923; // @[Mul.scala 207:34]
  wire  sum_1031 = sum_926 ^ sum_927; // @[Mul.scala 206:34]
  wire  cout_1031 = sum_926 & sum_927; // @[Mul.scala 207:34]
  wire  sum_1032 = cout_924 ^ cout_925; // @[Mul.scala 206:34]
  wire  cout_1032 = cout_924 & cout_925; // @[Mul.scala 207:34]
  wire  sum_1033 = sum_928 ^ sum_929; // @[Mul.scala 206:34]
  wire  cout_1033 = sum_928 & sum_929; // @[Mul.scala 207:34]
  wire  sum_1034 = cout_926 ^ cout_927; // @[Mul.scala 206:34]
  wire  cout_1034 = cout_926 & cout_927; // @[Mul.scala 207:34]
  wire  sum_1035 = sum_930 ^ sum_931; // @[Mul.scala 206:34]
  wire  cout_1035 = sum_930 & sum_931; // @[Mul.scala 207:34]
  wire  sum_1036 = cout_928 ^ cout_929; // @[Mul.scala 206:34]
  wire  cout_1036 = cout_928 & cout_929; // @[Mul.scala 207:34]
  wire  sum_1037 = sum_932 ^ sum_933; // @[Mul.scala 206:34]
  wire  cout_1037 = sum_932 & sum_933; // @[Mul.scala 207:34]
  wire  sum_1038 = cout_930 ^ cout_931; // @[Mul.scala 206:34]
  wire  cout_1038 = cout_930 & cout_931; // @[Mul.scala 207:34]
  wire  sum_1039 = sum_934 ^ sum_935; // @[Mul.scala 206:34]
  wire  cout_1039 = sum_934 & sum_935; // @[Mul.scala 207:34]
  wire  sum_1040 = cout_932 ^ cout_933; // @[Mul.scala 206:34]
  wire  cout_1040 = cout_932 & cout_933; // @[Mul.scala 207:34]
  wire  sum_1041 = sum_936 ^ sum_937; // @[Mul.scala 206:34]
  wire  cout_1041 = sum_936 & sum_937; // @[Mul.scala 207:34]
  wire  sum_1042 = cout_934 ^ cout_935; // @[Mul.scala 206:34]
  wire  cout_1042 = cout_934 & cout_935; // @[Mul.scala 207:34]
  wire  sum_1043 = sum_938 ^ sum_939; // @[Mul.scala 206:34]
  wire  cout_1043 = sum_938 & sum_939; // @[Mul.scala 207:34]
  wire  sum_1044 = cout_936 ^ cout_937; // @[Mul.scala 206:34]
  wire  cout_1044 = cout_936 & cout_937; // @[Mul.scala 207:34]
  wire  sum_1045 = sum_940 ^ sum_941; // @[Mul.scala 206:34]
  wire  cout_1045 = sum_940 & sum_941; // @[Mul.scala 207:34]
  wire  sum_1046 = cout_938 ^ cout_939; // @[Mul.scala 206:34]
  wire  cout_1046 = cout_938 & cout_939; // @[Mul.scala 207:34]
  wire  sum_1047 = sum_942 ^ sum_943; // @[Mul.scala 206:34]
  wire  cout_1047 = sum_942 & sum_943; // @[Mul.scala 207:34]
  wire  sum_1048 = cout_940 ^ cout_941; // @[Mul.scala 206:34]
  wire  cout_1048 = cout_940 & cout_941; // @[Mul.scala 207:34]
  wire  sum_1049 = sum_944 ^ sum_945; // @[Mul.scala 206:34]
  wire  cout_1049 = sum_944 & sum_945; // @[Mul.scala 207:34]
  wire  sum_1050 = cout_942 ^ cout_943; // @[Mul.scala 206:34]
  wire  cout_1050 = cout_942 & cout_943; // @[Mul.scala 207:34]
  wire  sum_1051 = sum_946 ^ sum_947; // @[Mul.scala 206:34]
  wire  cout_1051 = sum_946 & sum_947; // @[Mul.scala 207:34]
  wire  sum_1052 = cout_944 ^ cout_945; // @[Mul.scala 206:34]
  wire  cout_1052 = cout_944 & cout_945; // @[Mul.scala 207:34]
  wire  sum_1053 = sum_948 ^ sum_949; // @[Mul.scala 206:34]
  wire  cout_1053 = sum_948 & sum_949; // @[Mul.scala 207:34]
  wire  sum_1054 = cout_946 ^ cout_947; // @[Mul.scala 206:34]
  wire  cout_1054 = cout_946 & cout_947; // @[Mul.scala 207:34]
  wire  sum_1055 = sum_950 ^ sum_951; // @[Mul.scala 206:34]
  wire  cout_1055 = sum_950 & sum_951; // @[Mul.scala 207:34]
  wire  sum_1056 = cout_948 ^ cout_949; // @[Mul.scala 206:34]
  wire  cout_1056 = cout_948 & cout_949; // @[Mul.scala 207:34]
  wire  sum_1057 = sum_952 ^ sum_953; // @[Mul.scala 206:34]
  wire  cout_1057 = sum_952 & sum_953; // @[Mul.scala 207:34]
  wire  sum_1058 = cout_950 ^ cout_951; // @[Mul.scala 206:34]
  wire  cout_1058 = cout_950 & cout_951; // @[Mul.scala 207:34]
  wire  sum_1059 = sum_954 ^ sum_955; // @[Mul.scala 206:34]
  wire  cout_1059 = sum_954 & sum_955; // @[Mul.scala 207:34]
  wire  sum_1060 = cout_952 ^ cout_953; // @[Mul.scala 206:34]
  wire  cout_1060 = cout_952 & cout_953; // @[Mul.scala 207:34]
  wire  sum_1061 = sum_956 ^ sum_957; // @[Mul.scala 206:34]
  wire  cout_1061 = sum_956 & sum_957; // @[Mul.scala 207:34]
  wire  sum_1062 = cout_954 ^ cout_955; // @[Mul.scala 206:34]
  wire  cout_1062 = cout_954 & cout_955; // @[Mul.scala 207:34]
  wire  sum_1063 = sum_958 ^ sum_959; // @[Mul.scala 206:34]
  wire  cout_1063 = sum_958 & sum_959; // @[Mul.scala 207:34]
  wire  sum_1064 = cout_956 ^ cout_957; // @[Mul.scala 206:34]
  wire  cout_1064 = cout_956 & cout_957; // @[Mul.scala 207:34]
  wire  _sum_T_1685 = sum_960 ^ cout_958; // @[Mul.scala 191:34]
  wire  sum_1065 = sum_960 ^ cout_958 ^ cout_959; // @[Mul.scala 191:42]
  wire  cout_1065 = sum_960 & cout_958 | _sum_T_1685 & cout_959; // @[Mul.scala 192:44]
  wire  sum_1066 = sum_961 ^ cout_960; // @[Mul.scala 206:34]
  wire  cout_1066 = sum_961 & cout_960; // @[Mul.scala 207:34]
  wire  sum_1067 = sum_962 ^ cout_961; // @[Mul.scala 206:34]
  wire  cout_1067 = sum_962 & cout_961; // @[Mul.scala 207:34]
  wire  sum_1068 = sum_963 ^ cout_962; // @[Mul.scala 206:34]
  wire  cout_1068 = sum_963 & cout_962; // @[Mul.scala 207:34]
  wire  sum_1069 = sum_964 ^ cout_963; // @[Mul.scala 206:34]
  wire  cout_1069 = sum_964 & cout_963; // @[Mul.scala 207:34]
  wire  sum_1070 = sum_965 ^ cout_964; // @[Mul.scala 206:34]
  wire  sum_1083 = sum_978 ^ cout_977; // @[Mul.scala 206:34]
  wire  cout_1083 = sum_978 & cout_977; // @[Mul.scala 207:34]
  wire  sum_1084 = sum_979 ^ cout_978; // @[Mul.scala 206:34]
  wire  cout_1084 = sum_979 & cout_978; // @[Mul.scala 207:34]
  wire  sum_1085 = sum_980 ^ cout_979; // @[Mul.scala 206:34]
  wire  cout_1085 = sum_980 & cout_979; // @[Mul.scala 207:34]
  wire  _sum_T_1707 = sum_981 ^ sum_982; // @[Mul.scala 191:34]
  wire  sum_1086 = sum_981 ^ sum_982 ^ cout_980; // @[Mul.scala 191:42]
  wire  cout_1086 = sum_981 & sum_982 | _sum_T_1707 & cout_980; // @[Mul.scala 192:44]
  wire  sum_1087 = sum_983 ^ sum_984; // @[Mul.scala 206:34]
  wire  cout_1087 = sum_983 & sum_984; // @[Mul.scala 207:34]
  wire  sum_1088 = cout_981 ^ cout_982; // @[Mul.scala 206:34]
  wire  cout_1088 = cout_981 & cout_982; // @[Mul.scala 207:34]
  wire  sum_1089 = sum_985 ^ sum_986; // @[Mul.scala 206:34]
  wire  cout_1089 = sum_985 & sum_986; // @[Mul.scala 207:34]
  wire  sum_1090 = cout_983 ^ cout_984; // @[Mul.scala 206:34]
  wire  cout_1090 = cout_983 & cout_984; // @[Mul.scala 207:34]
  wire  sum_1091 = sum_987 ^ sum_988; // @[Mul.scala 206:34]
  wire  cout_1091 = sum_987 & sum_988; // @[Mul.scala 207:34]
  wire  sum_1092 = cout_985 ^ cout_986; // @[Mul.scala 206:34]
  wire  cout_1092 = cout_985 & cout_986; // @[Mul.scala 207:34]
  wire  sum_1093 = sum_989 ^ sum_990; // @[Mul.scala 206:34]
  wire  cout_1093 = sum_989 & sum_990; // @[Mul.scala 207:34]
  wire  sum_1094 = cout_987 ^ cout_988; // @[Mul.scala 206:34]
  wire  cout_1094 = cout_987 & cout_988; // @[Mul.scala 207:34]
  wire  sum_1095 = sum_991 ^ sum_992; // @[Mul.scala 206:34]
  wire  cout_1095 = sum_991 & sum_992; // @[Mul.scala 207:34]
  wire  sum_1096 = cout_989 ^ cout_990; // @[Mul.scala 206:34]
  wire  cout_1096 = cout_989 & cout_990; // @[Mul.scala 207:34]
  wire  sum_1097 = sum_993 ^ sum_994; // @[Mul.scala 206:34]
  wire  cout_1097 = sum_993 & sum_994; // @[Mul.scala 207:34]
  wire  sum_1098 = cout_991 ^ cout_992; // @[Mul.scala 206:34]
  wire  cout_1098 = cout_991 & cout_992; // @[Mul.scala 207:34]
  wire  sum_1099 = sum_995 ^ sum_996; // @[Mul.scala 206:34]
  wire  cout_1099 = sum_995 & sum_996; // @[Mul.scala 207:34]
  wire  sum_1100 = cout_993 ^ cout_994; // @[Mul.scala 206:34]
  wire  cout_1100 = cout_993 & cout_994; // @[Mul.scala 207:34]
  wire  sum_1101 = sum_997 ^ sum_998; // @[Mul.scala 206:34]
  wire  cout_1101 = sum_997 & sum_998; // @[Mul.scala 207:34]
  wire  sum_1102 = cout_995 ^ cout_996; // @[Mul.scala 206:34]
  wire  cout_1102 = cout_995 & cout_996; // @[Mul.scala 207:34]
  wire  sum_1103 = sum_999 ^ sum_1000; // @[Mul.scala 206:34]
  wire  cout_1103 = sum_999 & sum_1000; // @[Mul.scala 207:34]
  wire  sum_1104 = cout_997 ^ cout_998; // @[Mul.scala 206:34]
  wire  cout_1104 = cout_997 & cout_998; // @[Mul.scala 207:34]
  wire  sum_1105 = sum_1001 ^ sum_1002; // @[Mul.scala 206:34]
  wire  cout_1105 = sum_1001 & sum_1002; // @[Mul.scala 207:34]
  wire  sum_1106 = cout_999 ^ cout_1000; // @[Mul.scala 206:34]
  wire  cout_1106 = cout_999 & cout_1000; // @[Mul.scala 207:34]
  wire  sum_1107 = sum_1003 ^ sum_1004; // @[Mul.scala 206:34]
  wire  cout_1107 = sum_1003 & sum_1004; // @[Mul.scala 207:34]
  wire  sum_1108 = cout_1001 ^ cout_1002; // @[Mul.scala 206:34]
  wire  cout_1108 = cout_1001 & cout_1002; // @[Mul.scala 207:34]
  wire  sum_1109 = sum_1005 ^ sum_1006; // @[Mul.scala 206:34]
  wire  cout_1109 = sum_1005 & sum_1006; // @[Mul.scala 207:34]
  wire  sum_1110 = cout_1003 ^ cout_1004; // @[Mul.scala 206:34]
  wire  cout_1110 = cout_1003 & cout_1004; // @[Mul.scala 207:34]
  wire  sum_1111 = sum_1007 ^ sum_1008; // @[Mul.scala 206:34]
  wire  cout_1111 = sum_1007 & sum_1008; // @[Mul.scala 207:34]
  wire  sum_1112 = cout_1005 ^ cout_1006; // @[Mul.scala 206:34]
  wire  cout_1112 = cout_1005 & cout_1006; // @[Mul.scala 207:34]
  wire  sum_1113 = sum_1009 ^ sum_1010; // @[Mul.scala 206:34]
  wire  cout_1113 = sum_1009 & sum_1010; // @[Mul.scala 207:34]
  wire  sum_1114 = cout_1007 ^ cout_1008; // @[Mul.scala 206:34]
  wire  cout_1114 = cout_1007 & cout_1008; // @[Mul.scala 207:34]
  wire  sum_1115 = sum_1011 ^ sum_1012; // @[Mul.scala 206:34]
  wire  cout_1115 = sum_1011 & sum_1012; // @[Mul.scala 207:34]
  wire  sum_1116 = cout_1009 ^ cout_1010; // @[Mul.scala 206:34]
  wire  cout_1116 = cout_1009 & cout_1010; // @[Mul.scala 207:34]
  wire  sum_1117 = sum_1013 ^ sum_1014; // @[Mul.scala 206:34]
  wire  cout_1117 = sum_1013 & sum_1014; // @[Mul.scala 207:34]
  wire  sum_1118 = cout_1011 ^ cout_1012; // @[Mul.scala 206:34]
  wire  cout_1118 = cout_1011 & cout_1012; // @[Mul.scala 207:34]
  wire  sum_1119 = sum_1015 ^ sum_1016; // @[Mul.scala 206:34]
  wire  cout_1119 = sum_1015 & sum_1016; // @[Mul.scala 207:34]
  wire  sum_1120 = cout_1013 ^ cout_1014; // @[Mul.scala 206:34]
  wire  cout_1120 = cout_1013 & cout_1014; // @[Mul.scala 207:34]
  wire  sum_1121 = sum_1017 ^ sum_1018; // @[Mul.scala 206:34]
  wire  cout_1121 = sum_1017 & sum_1018; // @[Mul.scala 207:34]
  wire  sum_1122 = cout_1015 ^ cout_1016; // @[Mul.scala 206:34]
  wire  cout_1122 = cout_1015 & cout_1016; // @[Mul.scala 207:34]
  wire  sum_1123 = sum_1019 ^ sum_1020; // @[Mul.scala 206:34]
  wire  cout_1123 = sum_1019 & sum_1020; // @[Mul.scala 207:34]
  wire  sum_1124 = cout_1017 ^ cout_1018; // @[Mul.scala 206:34]
  wire  cout_1124 = cout_1017 & cout_1018; // @[Mul.scala 207:34]
  wire  sum_1125 = sum_1021 ^ sum_1022; // @[Mul.scala 206:34]
  wire  cout_1125 = sum_1021 & sum_1022; // @[Mul.scala 207:34]
  wire  sum_1126 = cout_1019 ^ cout_1020; // @[Mul.scala 206:34]
  wire  cout_1126 = cout_1019 & cout_1020; // @[Mul.scala 207:34]
  wire  sum_1127 = sum_1023 ^ sum_1024; // @[Mul.scala 206:34]
  wire  cout_1127 = sum_1023 & sum_1024; // @[Mul.scala 207:34]
  wire  sum_1128 = cout_1021 ^ cout_1022; // @[Mul.scala 206:34]
  wire  cout_1128 = cout_1021 & cout_1022; // @[Mul.scala 207:34]
  wire  sum_1129 = sum_1025 ^ sum_1026; // @[Mul.scala 206:34]
  wire  cout_1129 = sum_1025 & sum_1026; // @[Mul.scala 207:34]
  wire  sum_1130 = cout_1023 ^ cout_1024; // @[Mul.scala 206:34]
  wire  cout_1130 = cout_1023 & cout_1024; // @[Mul.scala 207:34]
  wire  sum_1131 = sum_1027 ^ sum_1028; // @[Mul.scala 206:34]
  wire  cout_1131 = sum_1027 & sum_1028; // @[Mul.scala 207:34]
  wire  sum_1132 = cout_1025 ^ cout_1026; // @[Mul.scala 206:34]
  wire  cout_1132 = cout_1025 & cout_1026; // @[Mul.scala 207:34]
  wire  sum_1133 = sum_1029 ^ sum_1030; // @[Mul.scala 206:34]
  wire  cout_1133 = sum_1029 & sum_1030; // @[Mul.scala 207:34]
  wire  sum_1134 = cout_1027 ^ cout_1028; // @[Mul.scala 206:34]
  wire  cout_1134 = cout_1027 & cout_1028; // @[Mul.scala 207:34]
  wire  sum_1135 = sum_1031 ^ sum_1032; // @[Mul.scala 206:34]
  wire  cout_1135 = sum_1031 & sum_1032; // @[Mul.scala 207:34]
  wire  sum_1136 = cout_1029 ^ cout_1030; // @[Mul.scala 206:34]
  wire  cout_1136 = cout_1029 & cout_1030; // @[Mul.scala 207:34]
  wire  sum_1137 = sum_1033 ^ sum_1034; // @[Mul.scala 206:34]
  wire  cout_1137 = sum_1033 & sum_1034; // @[Mul.scala 207:34]
  wire  sum_1138 = cout_1031 ^ cout_1032; // @[Mul.scala 206:34]
  wire  cout_1138 = cout_1031 & cout_1032; // @[Mul.scala 207:34]
  wire  sum_1139 = sum_1035 ^ sum_1036; // @[Mul.scala 206:34]
  wire  cout_1139 = sum_1035 & sum_1036; // @[Mul.scala 207:34]
  wire  sum_1140 = cout_1033 ^ cout_1034; // @[Mul.scala 206:34]
  wire  cout_1140 = cout_1033 & cout_1034; // @[Mul.scala 207:34]
  wire  sum_1141 = sum_1037 ^ sum_1038; // @[Mul.scala 206:34]
  wire  cout_1141 = sum_1037 & sum_1038; // @[Mul.scala 207:34]
  wire  sum_1142 = cout_1035 ^ cout_1036; // @[Mul.scala 206:34]
  wire  cout_1142 = cout_1035 & cout_1036; // @[Mul.scala 207:34]
  wire  sum_1143 = sum_1039 ^ sum_1040; // @[Mul.scala 206:34]
  wire  cout_1143 = sum_1039 & sum_1040; // @[Mul.scala 207:34]
  wire  sum_1144 = cout_1037 ^ cout_1038; // @[Mul.scala 206:34]
  wire  cout_1144 = cout_1037 & cout_1038; // @[Mul.scala 207:34]
  wire  sum_1145 = sum_1041 ^ sum_1042; // @[Mul.scala 206:34]
  wire  cout_1145 = sum_1041 & sum_1042; // @[Mul.scala 207:34]
  wire  sum_1146 = cout_1039 ^ cout_1040; // @[Mul.scala 206:34]
  wire  cout_1146 = cout_1039 & cout_1040; // @[Mul.scala 207:34]
  wire  sum_1147 = sum_1043 ^ sum_1044; // @[Mul.scala 206:34]
  wire  cout_1147 = sum_1043 & sum_1044; // @[Mul.scala 207:34]
  wire  sum_1148 = cout_1041 ^ cout_1042; // @[Mul.scala 206:34]
  wire  cout_1148 = cout_1041 & cout_1042; // @[Mul.scala 207:34]
  wire  sum_1149 = sum_1045 ^ sum_1046; // @[Mul.scala 206:34]
  wire  cout_1149 = sum_1045 & sum_1046; // @[Mul.scala 207:34]
  wire  sum_1150 = cout_1043 ^ cout_1044; // @[Mul.scala 206:34]
  wire  cout_1150 = cout_1043 & cout_1044; // @[Mul.scala 207:34]
  wire  sum_1151 = sum_1047 ^ sum_1048; // @[Mul.scala 206:34]
  wire  cout_1151 = sum_1047 & sum_1048; // @[Mul.scala 207:34]
  wire  sum_1152 = cout_1045 ^ cout_1046; // @[Mul.scala 206:34]
  wire  cout_1152 = cout_1045 & cout_1046; // @[Mul.scala 207:34]
  wire  sum_1153 = sum_1049 ^ sum_1050; // @[Mul.scala 206:34]
  wire  cout_1153 = sum_1049 & sum_1050; // @[Mul.scala 207:34]
  wire  sum_1154 = cout_1047 ^ cout_1048; // @[Mul.scala 206:34]
  wire  cout_1154 = cout_1047 & cout_1048; // @[Mul.scala 207:34]
  wire  sum_1155 = sum_1051 ^ sum_1052; // @[Mul.scala 206:34]
  wire  cout_1155 = sum_1051 & sum_1052; // @[Mul.scala 207:34]
  wire  sum_1156 = cout_1049 ^ cout_1050; // @[Mul.scala 206:34]
  wire  cout_1156 = cout_1049 & cout_1050; // @[Mul.scala 207:34]
  wire  sum_1157 = sum_1053 ^ sum_1054; // @[Mul.scala 206:34]
  wire  cout_1157 = sum_1053 & sum_1054; // @[Mul.scala 207:34]
  wire  sum_1158 = cout_1051 ^ cout_1052; // @[Mul.scala 206:34]
  wire  cout_1158 = cout_1051 & cout_1052; // @[Mul.scala 207:34]
  wire  sum_1159 = sum_1055 ^ sum_1056; // @[Mul.scala 206:34]
  wire  cout_1159 = sum_1055 & sum_1056; // @[Mul.scala 207:34]
  wire  sum_1160 = cout_1053 ^ cout_1054; // @[Mul.scala 206:34]
  wire  cout_1160 = cout_1053 & cout_1054; // @[Mul.scala 207:34]
  wire  sum_1161 = sum_1057 ^ sum_1058; // @[Mul.scala 206:34]
  wire  cout_1161 = sum_1057 & sum_1058; // @[Mul.scala 207:34]
  wire  sum_1162 = cout_1055 ^ cout_1056; // @[Mul.scala 206:34]
  wire  cout_1162 = cout_1055 & cout_1056; // @[Mul.scala 207:34]
  wire  sum_1163 = sum_1059 ^ sum_1060; // @[Mul.scala 206:34]
  wire  cout_1163 = sum_1059 & sum_1060; // @[Mul.scala 207:34]
  wire  sum_1164 = cout_1057 ^ cout_1058; // @[Mul.scala 206:34]
  wire  cout_1164 = cout_1057 & cout_1058; // @[Mul.scala 207:34]
  wire  sum_1165 = sum_1061 ^ sum_1062; // @[Mul.scala 206:34]
  wire  cout_1165 = sum_1061 & sum_1062; // @[Mul.scala 207:34]
  wire  sum_1166 = cout_1059 ^ cout_1060; // @[Mul.scala 206:34]
  wire  cout_1166 = cout_1059 & cout_1060; // @[Mul.scala 207:34]
  wire  sum_1167 = sum_1063 ^ sum_1064; // @[Mul.scala 206:34]
  wire  cout_1167 = sum_1063 & sum_1064; // @[Mul.scala 207:34]
  wire  sum_1168 = cout_1061 ^ cout_1062; // @[Mul.scala 206:34]
  wire  cout_1168 = cout_1061 & cout_1062; // @[Mul.scala 207:34]
  wire  _sum_T_1791 = sum_1065 ^ cout_1063; // @[Mul.scala 191:34]
  wire  sum_1169 = sum_1065 ^ cout_1063 ^ cout_1064; // @[Mul.scala 191:42]
  wire  cout_1169 = sum_1065 & cout_1063 | _sum_T_1791 & cout_1064; // @[Mul.scala 192:44]
  wire  sum_1170 = sum_1066 ^ cout_1065; // @[Mul.scala 206:34]
  wire  cout_1170 = sum_1066 & cout_1065; // @[Mul.scala 207:34]
  wire  sum_1171 = sum_1067 ^ cout_1066; // @[Mul.scala 206:34]
  wire  cout_1171 = sum_1067 & cout_1066; // @[Mul.scala 207:34]
  wire  sum_1172 = sum_1068 ^ cout_1067; // @[Mul.scala 206:34]
  wire  cout_1172 = sum_1068 & cout_1067; // @[Mul.scala 207:34]
  wire  sum_1173 = sum_1069 ^ cout_1068; // @[Mul.scala 206:34]
  wire  cout_1173 = sum_1069 & cout_1068; // @[Mul.scala 207:34]
  wire  sum_1174 = sum_1070 ^ cout_1069; // @[Mul.scala 206:34]
  wire  sum_1188 = sum_1084 ^ cout_1083; // @[Mul.scala 206:34]
  wire  cout_1188 = sum_1084 & cout_1083; // @[Mul.scala 207:34]
  wire  sum_1189 = sum_1085 ^ cout_1084; // @[Mul.scala 206:34]
  wire  cout_1189 = sum_1085 & cout_1084; // @[Mul.scala 207:34]
  wire  sum_1190 = sum_1086 ^ cout_1085; // @[Mul.scala 206:34]
  wire  cout_1190 = sum_1086 & cout_1085; // @[Mul.scala 207:34]
  wire  _sum_T_1814 = sum_1087 ^ sum_1088; // @[Mul.scala 191:34]
  wire  sum_1191 = sum_1087 ^ sum_1088 ^ cout_1086; // @[Mul.scala 191:42]
  wire  cout_1191 = sum_1087 & sum_1088 | _sum_T_1814 & cout_1086; // @[Mul.scala 192:44]
  wire  sum_1192 = sum_1089 ^ sum_1090; // @[Mul.scala 206:34]
  wire  cout_1192 = sum_1089 & sum_1090; // @[Mul.scala 207:34]
  wire  sum_1193 = cout_1087 ^ cout_1088; // @[Mul.scala 206:34]
  wire  cout_1193 = cout_1087 & cout_1088; // @[Mul.scala 207:34]
  wire  sum_1194 = sum_1091 ^ sum_1092; // @[Mul.scala 206:34]
  wire  cout_1194 = sum_1091 & sum_1092; // @[Mul.scala 207:34]
  wire  sum_1195 = cout_1089 ^ cout_1090; // @[Mul.scala 206:34]
  wire  cout_1195 = cout_1089 & cout_1090; // @[Mul.scala 207:34]
  wire  sum_1196 = sum_1093 ^ sum_1094; // @[Mul.scala 206:34]
  wire  cout_1196 = sum_1093 & sum_1094; // @[Mul.scala 207:34]
  wire  sum_1197 = cout_1091 ^ cout_1092; // @[Mul.scala 206:34]
  wire  cout_1197 = cout_1091 & cout_1092; // @[Mul.scala 207:34]
  wire  sum_1198 = sum_1095 ^ sum_1096; // @[Mul.scala 206:34]
  wire  cout_1198 = sum_1095 & sum_1096; // @[Mul.scala 207:34]
  wire  sum_1199 = cout_1093 ^ cout_1094; // @[Mul.scala 206:34]
  wire  cout_1199 = cout_1093 & cout_1094; // @[Mul.scala 207:34]
  wire  sum_1200 = sum_1097 ^ sum_1098; // @[Mul.scala 206:34]
  wire  cout_1200 = sum_1097 & sum_1098; // @[Mul.scala 207:34]
  wire  sum_1201 = cout_1095 ^ cout_1096; // @[Mul.scala 206:34]
  wire  cout_1201 = cout_1095 & cout_1096; // @[Mul.scala 207:34]
  wire  sum_1202 = sum_1099 ^ sum_1100; // @[Mul.scala 206:34]
  wire  cout_1202 = sum_1099 & sum_1100; // @[Mul.scala 207:34]
  wire  sum_1203 = cout_1097 ^ cout_1098; // @[Mul.scala 206:34]
  wire  cout_1203 = cout_1097 & cout_1098; // @[Mul.scala 207:34]
  wire  sum_1204 = sum_1101 ^ sum_1102; // @[Mul.scala 206:34]
  wire  cout_1204 = sum_1101 & sum_1102; // @[Mul.scala 207:34]
  wire  sum_1205 = cout_1099 ^ cout_1100; // @[Mul.scala 206:34]
  wire  cout_1205 = cout_1099 & cout_1100; // @[Mul.scala 207:34]
  wire  sum_1206 = sum_1103 ^ sum_1104; // @[Mul.scala 206:34]
  wire  cout_1206 = sum_1103 & sum_1104; // @[Mul.scala 207:34]
  wire  sum_1207 = cout_1101 ^ cout_1102; // @[Mul.scala 206:34]
  wire  cout_1207 = cout_1101 & cout_1102; // @[Mul.scala 207:34]
  wire  sum_1208 = sum_1105 ^ sum_1106; // @[Mul.scala 206:34]
  wire  cout_1208 = sum_1105 & sum_1106; // @[Mul.scala 207:34]
  wire  sum_1209 = cout_1103 ^ cout_1104; // @[Mul.scala 206:34]
  wire  cout_1209 = cout_1103 & cout_1104; // @[Mul.scala 207:34]
  wire  sum_1210 = sum_1107 ^ sum_1108; // @[Mul.scala 206:34]
  wire  cout_1210 = sum_1107 & sum_1108; // @[Mul.scala 207:34]
  wire  sum_1211 = cout_1105 ^ cout_1106; // @[Mul.scala 206:34]
  wire  cout_1211 = cout_1105 & cout_1106; // @[Mul.scala 207:34]
  wire  sum_1212 = sum_1109 ^ sum_1110; // @[Mul.scala 206:34]
  wire  cout_1212 = sum_1109 & sum_1110; // @[Mul.scala 207:34]
  wire  sum_1213 = cout_1107 ^ cout_1108; // @[Mul.scala 206:34]
  wire  cout_1213 = cout_1107 & cout_1108; // @[Mul.scala 207:34]
  wire  sum_1214 = sum_1111 ^ sum_1112; // @[Mul.scala 206:34]
  wire  cout_1214 = sum_1111 & sum_1112; // @[Mul.scala 207:34]
  wire  sum_1215 = cout_1109 ^ cout_1110; // @[Mul.scala 206:34]
  wire  cout_1215 = cout_1109 & cout_1110; // @[Mul.scala 207:34]
  wire  sum_1216 = sum_1113 ^ sum_1114; // @[Mul.scala 206:34]
  wire  cout_1216 = sum_1113 & sum_1114; // @[Mul.scala 207:34]
  wire  sum_1217 = cout_1111 ^ cout_1112; // @[Mul.scala 206:34]
  wire  cout_1217 = cout_1111 & cout_1112; // @[Mul.scala 207:34]
  wire  sum_1218 = sum_1115 ^ sum_1116; // @[Mul.scala 206:34]
  wire  cout_1218 = sum_1115 & sum_1116; // @[Mul.scala 207:34]
  wire  sum_1219 = cout_1113 ^ cout_1114; // @[Mul.scala 206:34]
  wire  cout_1219 = cout_1113 & cout_1114; // @[Mul.scala 207:34]
  wire  sum_1220 = sum_1117 ^ sum_1118; // @[Mul.scala 206:34]
  wire  cout_1220 = sum_1117 & sum_1118; // @[Mul.scala 207:34]
  wire  sum_1221 = cout_1115 ^ cout_1116; // @[Mul.scala 206:34]
  wire  cout_1221 = cout_1115 & cout_1116; // @[Mul.scala 207:34]
  wire  sum_1222 = sum_1119 ^ sum_1120; // @[Mul.scala 206:34]
  wire  cout_1222 = sum_1119 & sum_1120; // @[Mul.scala 207:34]
  wire  sum_1223 = cout_1117 ^ cout_1118; // @[Mul.scala 206:34]
  wire  cout_1223 = cout_1117 & cout_1118; // @[Mul.scala 207:34]
  wire  sum_1224 = sum_1121 ^ sum_1122; // @[Mul.scala 206:34]
  wire  cout_1224 = sum_1121 & sum_1122; // @[Mul.scala 207:34]
  wire  sum_1225 = cout_1119 ^ cout_1120; // @[Mul.scala 206:34]
  wire  cout_1225 = cout_1119 & cout_1120; // @[Mul.scala 207:34]
  wire  sum_1226 = sum_1123 ^ sum_1124; // @[Mul.scala 206:34]
  wire  cout_1226 = sum_1123 & sum_1124; // @[Mul.scala 207:34]
  wire  sum_1227 = cout_1121 ^ cout_1122; // @[Mul.scala 206:34]
  wire  cout_1227 = cout_1121 & cout_1122; // @[Mul.scala 207:34]
  wire  sum_1228 = sum_1125 ^ sum_1126; // @[Mul.scala 206:34]
  wire  cout_1228 = sum_1125 & sum_1126; // @[Mul.scala 207:34]
  wire  sum_1229 = cout_1123 ^ cout_1124; // @[Mul.scala 206:34]
  wire  cout_1229 = cout_1123 & cout_1124; // @[Mul.scala 207:34]
  wire  sum_1230 = sum_1127 ^ sum_1128; // @[Mul.scala 206:34]
  wire  cout_1230 = sum_1127 & sum_1128; // @[Mul.scala 207:34]
  wire  sum_1231 = cout_1125 ^ cout_1126; // @[Mul.scala 206:34]
  wire  cout_1231 = cout_1125 & cout_1126; // @[Mul.scala 207:34]
  wire  sum_1232 = sum_1129 ^ sum_1130; // @[Mul.scala 206:34]
  wire  cout_1232 = sum_1129 & sum_1130; // @[Mul.scala 207:34]
  wire  sum_1233 = cout_1127 ^ cout_1128; // @[Mul.scala 206:34]
  wire  cout_1233 = cout_1127 & cout_1128; // @[Mul.scala 207:34]
  wire  sum_1234 = sum_1131 ^ sum_1132; // @[Mul.scala 206:34]
  wire  cout_1234 = sum_1131 & sum_1132; // @[Mul.scala 207:34]
  wire  sum_1235 = cout_1129 ^ cout_1130; // @[Mul.scala 206:34]
  wire  cout_1235 = cout_1129 & cout_1130; // @[Mul.scala 207:34]
  wire  sum_1236 = sum_1133 ^ sum_1134; // @[Mul.scala 206:34]
  wire  cout_1236 = sum_1133 & sum_1134; // @[Mul.scala 207:34]
  wire  sum_1237 = cout_1131 ^ cout_1132; // @[Mul.scala 206:34]
  wire  cout_1237 = cout_1131 & cout_1132; // @[Mul.scala 207:34]
  wire  sum_1238 = sum_1135 ^ sum_1136; // @[Mul.scala 206:34]
  wire  cout_1238 = sum_1135 & sum_1136; // @[Mul.scala 207:34]
  wire  sum_1239 = cout_1133 ^ cout_1134; // @[Mul.scala 206:34]
  wire  cout_1239 = cout_1133 & cout_1134; // @[Mul.scala 207:34]
  wire  sum_1240 = sum_1137 ^ sum_1138; // @[Mul.scala 206:34]
  wire  cout_1240 = sum_1137 & sum_1138; // @[Mul.scala 207:34]
  wire  sum_1241 = cout_1135 ^ cout_1136; // @[Mul.scala 206:34]
  wire  cout_1241 = cout_1135 & cout_1136; // @[Mul.scala 207:34]
  wire  sum_1242 = sum_1139 ^ sum_1140; // @[Mul.scala 206:34]
  wire  cout_1242 = sum_1139 & sum_1140; // @[Mul.scala 207:34]
  wire  sum_1243 = cout_1137 ^ cout_1138; // @[Mul.scala 206:34]
  wire  cout_1243 = cout_1137 & cout_1138; // @[Mul.scala 207:34]
  wire  sum_1244 = sum_1141 ^ sum_1142; // @[Mul.scala 206:34]
  wire  cout_1244 = sum_1141 & sum_1142; // @[Mul.scala 207:34]
  wire  sum_1245 = cout_1139 ^ cout_1140; // @[Mul.scala 206:34]
  wire  cout_1245 = cout_1139 & cout_1140; // @[Mul.scala 207:34]
  wire  sum_1246 = sum_1143 ^ sum_1144; // @[Mul.scala 206:34]
  wire  cout_1246 = sum_1143 & sum_1144; // @[Mul.scala 207:34]
  wire  sum_1247 = cout_1141 ^ cout_1142; // @[Mul.scala 206:34]
  wire  cout_1247 = cout_1141 & cout_1142; // @[Mul.scala 207:34]
  wire  sum_1248 = sum_1145 ^ sum_1146; // @[Mul.scala 206:34]
  wire  cout_1248 = sum_1145 & sum_1146; // @[Mul.scala 207:34]
  wire  sum_1249 = cout_1143 ^ cout_1144; // @[Mul.scala 206:34]
  wire  cout_1249 = cout_1143 & cout_1144; // @[Mul.scala 207:34]
  wire  sum_1250 = sum_1147 ^ sum_1148; // @[Mul.scala 206:34]
  wire  cout_1250 = sum_1147 & sum_1148; // @[Mul.scala 207:34]
  wire  sum_1251 = cout_1145 ^ cout_1146; // @[Mul.scala 206:34]
  wire  cout_1251 = cout_1145 & cout_1146; // @[Mul.scala 207:34]
  wire  sum_1252 = sum_1149 ^ sum_1150; // @[Mul.scala 206:34]
  wire  cout_1252 = sum_1149 & sum_1150; // @[Mul.scala 207:34]
  wire  sum_1253 = cout_1147 ^ cout_1148; // @[Mul.scala 206:34]
  wire  cout_1253 = cout_1147 & cout_1148; // @[Mul.scala 207:34]
  wire  sum_1254 = sum_1151 ^ sum_1152; // @[Mul.scala 206:34]
  wire  cout_1254 = sum_1151 & sum_1152; // @[Mul.scala 207:34]
  wire  sum_1255 = cout_1149 ^ cout_1150; // @[Mul.scala 206:34]
  wire  cout_1255 = cout_1149 & cout_1150; // @[Mul.scala 207:34]
  wire  sum_1256 = sum_1153 ^ sum_1154; // @[Mul.scala 206:34]
  wire  cout_1256 = sum_1153 & sum_1154; // @[Mul.scala 207:34]
  wire  sum_1257 = cout_1151 ^ cout_1152; // @[Mul.scala 206:34]
  wire  cout_1257 = cout_1151 & cout_1152; // @[Mul.scala 207:34]
  wire  sum_1258 = sum_1155 ^ sum_1156; // @[Mul.scala 206:34]
  wire  cout_1258 = sum_1155 & sum_1156; // @[Mul.scala 207:34]
  wire  sum_1259 = cout_1153 ^ cout_1154; // @[Mul.scala 206:34]
  wire  cout_1259 = cout_1153 & cout_1154; // @[Mul.scala 207:34]
  wire  sum_1260 = sum_1157 ^ sum_1158; // @[Mul.scala 206:34]
  wire  cout_1260 = sum_1157 & sum_1158; // @[Mul.scala 207:34]
  wire  sum_1261 = cout_1155 ^ cout_1156; // @[Mul.scala 206:34]
  wire  cout_1261 = cout_1155 & cout_1156; // @[Mul.scala 207:34]
  wire  sum_1262 = sum_1159 ^ sum_1160; // @[Mul.scala 206:34]
  wire  cout_1262 = sum_1159 & sum_1160; // @[Mul.scala 207:34]
  wire  sum_1263 = cout_1157 ^ cout_1158; // @[Mul.scala 206:34]
  wire  cout_1263 = cout_1157 & cout_1158; // @[Mul.scala 207:34]
  wire  sum_1264 = sum_1161 ^ sum_1162; // @[Mul.scala 206:34]
  wire  cout_1264 = sum_1161 & sum_1162; // @[Mul.scala 207:34]
  wire  sum_1265 = cout_1159 ^ cout_1160; // @[Mul.scala 206:34]
  wire  cout_1265 = cout_1159 & cout_1160; // @[Mul.scala 207:34]
  wire  sum_1266 = sum_1163 ^ sum_1164; // @[Mul.scala 206:34]
  wire  cout_1266 = sum_1163 & sum_1164; // @[Mul.scala 207:34]
  wire  sum_1267 = cout_1161 ^ cout_1162; // @[Mul.scala 206:34]
  wire  cout_1267 = cout_1161 & cout_1162; // @[Mul.scala 207:34]
  wire  sum_1268 = sum_1165 ^ sum_1166; // @[Mul.scala 206:34]
  wire  cout_1268 = sum_1165 & sum_1166; // @[Mul.scala 207:34]
  wire  sum_1269 = cout_1163 ^ cout_1164; // @[Mul.scala 206:34]
  wire  cout_1269 = cout_1163 & cout_1164; // @[Mul.scala 207:34]
  wire  sum_1270 = sum_1167 ^ sum_1168; // @[Mul.scala 206:34]
  wire  cout_1270 = sum_1167 & sum_1168; // @[Mul.scala 207:34]
  wire  sum_1271 = cout_1165 ^ cout_1166; // @[Mul.scala 206:34]
  wire  cout_1271 = cout_1165 & cout_1166; // @[Mul.scala 207:34]
  wire  _sum_T_1896 = sum_1169 ^ cout_1167; // @[Mul.scala 191:34]
  wire  sum_1272 = sum_1169 ^ cout_1167 ^ cout_1168; // @[Mul.scala 191:42]
  wire  cout_1272 = sum_1169 & cout_1167 | _sum_T_1896 & cout_1168; // @[Mul.scala 192:44]
  wire  sum_1273 = sum_1170 ^ cout_1169; // @[Mul.scala 206:34]
  wire  cout_1273 = sum_1170 & cout_1169; // @[Mul.scala 207:34]
  wire  sum_1274 = sum_1171 ^ cout_1170; // @[Mul.scala 206:34]
  wire  cout_1274 = sum_1171 & cout_1170; // @[Mul.scala 207:34]
  wire  sum_1275 = sum_1172 ^ cout_1171; // @[Mul.scala 206:34]
  wire  cout_1275 = sum_1172 & cout_1171; // @[Mul.scala 207:34]
  wire  sum_1276 = sum_1173 ^ cout_1172; // @[Mul.scala 206:34]
  wire  cout_1276 = sum_1173 & cout_1172; // @[Mul.scala 207:34]
  wire  sum_1277 = sum_1174 ^ cout_1173; // @[Mul.scala 206:34]
  wire  sum_1292 = sum_1189 ^ cout_1188; // @[Mul.scala 206:34]
  wire  cout_1292 = sum_1189 & cout_1188; // @[Mul.scala 207:34]
  wire  sum_1293 = sum_1190 ^ cout_1189; // @[Mul.scala 206:34]
  wire  cout_1293 = sum_1190 & cout_1189; // @[Mul.scala 207:34]
  wire  sum_1294 = sum_1191 ^ cout_1190; // @[Mul.scala 206:34]
  wire  cout_1294 = sum_1191 & cout_1190; // @[Mul.scala 207:34]
  wire  _sum_T_1920 = sum_1192 ^ sum_1193; // @[Mul.scala 191:34]
  wire  sum_1295 = sum_1192 ^ sum_1193 ^ cout_1191; // @[Mul.scala 191:42]
  wire  cout_1295 = sum_1192 & sum_1193 | _sum_T_1920 & cout_1191; // @[Mul.scala 192:44]
  wire  sum_1296 = sum_1194 ^ sum_1195; // @[Mul.scala 206:34]
  wire  cout_1296 = sum_1194 & sum_1195; // @[Mul.scala 207:34]
  wire  sum_1297 = cout_1192 ^ cout_1193; // @[Mul.scala 206:34]
  wire  cout_1297 = cout_1192 & cout_1193; // @[Mul.scala 207:34]
  wire  sum_1298 = sum_1196 ^ sum_1197; // @[Mul.scala 206:34]
  wire  cout_1298 = sum_1196 & sum_1197; // @[Mul.scala 207:34]
  wire  sum_1299 = cout_1194 ^ cout_1195; // @[Mul.scala 206:34]
  wire  cout_1299 = cout_1194 & cout_1195; // @[Mul.scala 207:34]
  wire  sum_1300 = sum_1198 ^ sum_1199; // @[Mul.scala 206:34]
  wire  cout_1300 = sum_1198 & sum_1199; // @[Mul.scala 207:34]
  wire  sum_1301 = cout_1196 ^ cout_1197; // @[Mul.scala 206:34]
  wire  cout_1301 = cout_1196 & cout_1197; // @[Mul.scala 207:34]
  wire  sum_1302 = sum_1200 ^ sum_1201; // @[Mul.scala 206:34]
  wire  cout_1302 = sum_1200 & sum_1201; // @[Mul.scala 207:34]
  wire  sum_1303 = cout_1198 ^ cout_1199; // @[Mul.scala 206:34]
  wire  cout_1303 = cout_1198 & cout_1199; // @[Mul.scala 207:34]
  wire  sum_1304 = sum_1202 ^ sum_1203; // @[Mul.scala 206:34]
  wire  cout_1304 = sum_1202 & sum_1203; // @[Mul.scala 207:34]
  wire  sum_1305 = cout_1200 ^ cout_1201; // @[Mul.scala 206:34]
  wire  cout_1305 = cout_1200 & cout_1201; // @[Mul.scala 207:34]
  wire  sum_1306 = sum_1204 ^ sum_1205; // @[Mul.scala 206:34]
  wire  cout_1306 = sum_1204 & sum_1205; // @[Mul.scala 207:34]
  wire  sum_1307 = cout_1202 ^ cout_1203; // @[Mul.scala 206:34]
  wire  cout_1307 = cout_1202 & cout_1203; // @[Mul.scala 207:34]
  wire  sum_1308 = sum_1206 ^ sum_1207; // @[Mul.scala 206:34]
  wire  cout_1308 = sum_1206 & sum_1207; // @[Mul.scala 207:34]
  wire  sum_1309 = cout_1204 ^ cout_1205; // @[Mul.scala 206:34]
  wire  cout_1309 = cout_1204 & cout_1205; // @[Mul.scala 207:34]
  wire  sum_1310 = sum_1208 ^ sum_1209; // @[Mul.scala 206:34]
  wire  cout_1310 = sum_1208 & sum_1209; // @[Mul.scala 207:34]
  wire  sum_1311 = cout_1206 ^ cout_1207; // @[Mul.scala 206:34]
  wire  cout_1311 = cout_1206 & cout_1207; // @[Mul.scala 207:34]
  wire  sum_1312 = sum_1210 ^ sum_1211; // @[Mul.scala 206:34]
  wire  cout_1312 = sum_1210 & sum_1211; // @[Mul.scala 207:34]
  wire  sum_1313 = cout_1208 ^ cout_1209; // @[Mul.scala 206:34]
  wire  cout_1313 = cout_1208 & cout_1209; // @[Mul.scala 207:34]
  wire  sum_1314 = sum_1212 ^ sum_1213; // @[Mul.scala 206:34]
  wire  cout_1314 = sum_1212 & sum_1213; // @[Mul.scala 207:34]
  wire  sum_1315 = cout_1210 ^ cout_1211; // @[Mul.scala 206:34]
  wire  cout_1315 = cout_1210 & cout_1211; // @[Mul.scala 207:34]
  wire  sum_1316 = sum_1214 ^ sum_1215; // @[Mul.scala 206:34]
  wire  cout_1316 = sum_1214 & sum_1215; // @[Mul.scala 207:34]
  wire  sum_1317 = cout_1212 ^ cout_1213; // @[Mul.scala 206:34]
  wire  cout_1317 = cout_1212 & cout_1213; // @[Mul.scala 207:34]
  wire  sum_1318 = sum_1216 ^ sum_1217; // @[Mul.scala 206:34]
  wire  cout_1318 = sum_1216 & sum_1217; // @[Mul.scala 207:34]
  wire  sum_1319 = cout_1214 ^ cout_1215; // @[Mul.scala 206:34]
  wire  cout_1319 = cout_1214 & cout_1215; // @[Mul.scala 207:34]
  wire  sum_1320 = sum_1218 ^ sum_1219; // @[Mul.scala 206:34]
  wire  cout_1320 = sum_1218 & sum_1219; // @[Mul.scala 207:34]
  wire  sum_1321 = cout_1216 ^ cout_1217; // @[Mul.scala 206:34]
  wire  cout_1321 = cout_1216 & cout_1217; // @[Mul.scala 207:34]
  wire  sum_1322 = sum_1220 ^ sum_1221; // @[Mul.scala 206:34]
  wire  cout_1322 = sum_1220 & sum_1221; // @[Mul.scala 207:34]
  wire  sum_1323 = cout_1218 ^ cout_1219; // @[Mul.scala 206:34]
  wire  cout_1323 = cout_1218 & cout_1219; // @[Mul.scala 207:34]
  wire  sum_1324 = sum_1222 ^ sum_1223; // @[Mul.scala 206:34]
  wire  cout_1324 = sum_1222 & sum_1223; // @[Mul.scala 207:34]
  wire  sum_1325 = cout_1220 ^ cout_1221; // @[Mul.scala 206:34]
  wire  cout_1325 = cout_1220 & cout_1221; // @[Mul.scala 207:34]
  wire  sum_1326 = sum_1224 ^ sum_1225; // @[Mul.scala 206:34]
  wire  cout_1326 = sum_1224 & sum_1225; // @[Mul.scala 207:34]
  wire  sum_1327 = cout_1222 ^ cout_1223; // @[Mul.scala 206:34]
  wire  cout_1327 = cout_1222 & cout_1223; // @[Mul.scala 207:34]
  wire  sum_1328 = sum_1226 ^ sum_1227; // @[Mul.scala 206:34]
  wire  cout_1328 = sum_1226 & sum_1227; // @[Mul.scala 207:34]
  wire  sum_1329 = cout_1224 ^ cout_1225; // @[Mul.scala 206:34]
  wire  cout_1329 = cout_1224 & cout_1225; // @[Mul.scala 207:34]
  wire  sum_1330 = sum_1228 ^ sum_1229; // @[Mul.scala 206:34]
  wire  cout_1330 = sum_1228 & sum_1229; // @[Mul.scala 207:34]
  wire  sum_1331 = cout_1226 ^ cout_1227; // @[Mul.scala 206:34]
  wire  cout_1331 = cout_1226 & cout_1227; // @[Mul.scala 207:34]
  wire  sum_1332 = sum_1230 ^ sum_1231; // @[Mul.scala 206:34]
  wire  cout_1332 = sum_1230 & sum_1231; // @[Mul.scala 207:34]
  wire  sum_1333 = cout_1228 ^ cout_1229; // @[Mul.scala 206:34]
  wire  cout_1333 = cout_1228 & cout_1229; // @[Mul.scala 207:34]
  wire  sum_1334 = sum_1232 ^ sum_1233; // @[Mul.scala 206:34]
  wire  cout_1334 = sum_1232 & sum_1233; // @[Mul.scala 207:34]
  wire  sum_1335 = cout_1230 ^ cout_1231; // @[Mul.scala 206:34]
  wire  cout_1335 = cout_1230 & cout_1231; // @[Mul.scala 207:34]
  wire  sum_1336 = sum_1234 ^ sum_1235; // @[Mul.scala 206:34]
  wire  cout_1336 = sum_1234 & sum_1235; // @[Mul.scala 207:34]
  wire  sum_1337 = cout_1232 ^ cout_1233; // @[Mul.scala 206:34]
  wire  cout_1337 = cout_1232 & cout_1233; // @[Mul.scala 207:34]
  wire  sum_1338 = sum_1236 ^ sum_1237; // @[Mul.scala 206:34]
  wire  cout_1338 = sum_1236 & sum_1237; // @[Mul.scala 207:34]
  wire  sum_1339 = cout_1234 ^ cout_1235; // @[Mul.scala 206:34]
  wire  cout_1339 = cout_1234 & cout_1235; // @[Mul.scala 207:34]
  wire  sum_1340 = sum_1238 ^ sum_1239; // @[Mul.scala 206:34]
  wire  cout_1340 = sum_1238 & sum_1239; // @[Mul.scala 207:34]
  wire  sum_1341 = cout_1236 ^ cout_1237; // @[Mul.scala 206:34]
  wire  cout_1341 = cout_1236 & cout_1237; // @[Mul.scala 207:34]
  wire  sum_1342 = sum_1240 ^ sum_1241; // @[Mul.scala 206:34]
  wire  cout_1342 = sum_1240 & sum_1241; // @[Mul.scala 207:34]
  wire  sum_1343 = cout_1238 ^ cout_1239; // @[Mul.scala 206:34]
  wire  cout_1343 = cout_1238 & cout_1239; // @[Mul.scala 207:34]
  wire  sum_1344 = sum_1242 ^ sum_1243; // @[Mul.scala 206:34]
  wire  cout_1344 = sum_1242 & sum_1243; // @[Mul.scala 207:34]
  wire  sum_1345 = cout_1240 ^ cout_1241; // @[Mul.scala 206:34]
  wire  cout_1345 = cout_1240 & cout_1241; // @[Mul.scala 207:34]
  wire  sum_1346 = sum_1244 ^ sum_1245; // @[Mul.scala 206:34]
  wire  cout_1346 = sum_1244 & sum_1245; // @[Mul.scala 207:34]
  wire  sum_1347 = cout_1242 ^ cout_1243; // @[Mul.scala 206:34]
  wire  cout_1347 = cout_1242 & cout_1243; // @[Mul.scala 207:34]
  wire  sum_1348 = sum_1246 ^ sum_1247; // @[Mul.scala 206:34]
  wire  cout_1348 = sum_1246 & sum_1247; // @[Mul.scala 207:34]
  wire  sum_1349 = cout_1244 ^ cout_1245; // @[Mul.scala 206:34]
  wire  cout_1349 = cout_1244 & cout_1245; // @[Mul.scala 207:34]
  wire  sum_1350 = sum_1248 ^ sum_1249; // @[Mul.scala 206:34]
  wire  cout_1350 = sum_1248 & sum_1249; // @[Mul.scala 207:34]
  wire  sum_1351 = cout_1246 ^ cout_1247; // @[Mul.scala 206:34]
  wire  cout_1351 = cout_1246 & cout_1247; // @[Mul.scala 207:34]
  wire  sum_1352 = sum_1250 ^ sum_1251; // @[Mul.scala 206:34]
  wire  cout_1352 = sum_1250 & sum_1251; // @[Mul.scala 207:34]
  wire  sum_1353 = cout_1248 ^ cout_1249; // @[Mul.scala 206:34]
  wire  cout_1353 = cout_1248 & cout_1249; // @[Mul.scala 207:34]
  wire  sum_1354 = sum_1252 ^ sum_1253; // @[Mul.scala 206:34]
  wire  cout_1354 = sum_1252 & sum_1253; // @[Mul.scala 207:34]
  wire  sum_1355 = cout_1250 ^ cout_1251; // @[Mul.scala 206:34]
  wire  cout_1355 = cout_1250 & cout_1251; // @[Mul.scala 207:34]
  wire  sum_1356 = sum_1254 ^ sum_1255; // @[Mul.scala 206:34]
  wire  cout_1356 = sum_1254 & sum_1255; // @[Mul.scala 207:34]
  wire  sum_1357 = cout_1252 ^ cout_1253; // @[Mul.scala 206:34]
  wire  cout_1357 = cout_1252 & cout_1253; // @[Mul.scala 207:34]
  wire  sum_1358 = sum_1256 ^ sum_1257; // @[Mul.scala 206:34]
  wire  cout_1358 = sum_1256 & sum_1257; // @[Mul.scala 207:34]
  wire  sum_1359 = cout_1254 ^ cout_1255; // @[Mul.scala 206:34]
  wire  cout_1359 = cout_1254 & cout_1255; // @[Mul.scala 207:34]
  wire  sum_1360 = sum_1258 ^ sum_1259; // @[Mul.scala 206:34]
  wire  cout_1360 = sum_1258 & sum_1259; // @[Mul.scala 207:34]
  wire  sum_1361 = cout_1256 ^ cout_1257; // @[Mul.scala 206:34]
  wire  cout_1361 = cout_1256 & cout_1257; // @[Mul.scala 207:34]
  wire  sum_1362 = sum_1260 ^ sum_1261; // @[Mul.scala 206:34]
  wire  cout_1362 = sum_1260 & sum_1261; // @[Mul.scala 207:34]
  wire  sum_1363 = cout_1258 ^ cout_1259; // @[Mul.scala 206:34]
  wire  cout_1363 = cout_1258 & cout_1259; // @[Mul.scala 207:34]
  wire  sum_1364 = sum_1262 ^ sum_1263; // @[Mul.scala 206:34]
  wire  cout_1364 = sum_1262 & sum_1263; // @[Mul.scala 207:34]
  wire  sum_1365 = cout_1260 ^ cout_1261; // @[Mul.scala 206:34]
  wire  cout_1365 = cout_1260 & cout_1261; // @[Mul.scala 207:34]
  wire  sum_1366 = sum_1264 ^ sum_1265; // @[Mul.scala 206:34]
  wire  cout_1366 = sum_1264 & sum_1265; // @[Mul.scala 207:34]
  wire  sum_1367 = cout_1262 ^ cout_1263; // @[Mul.scala 206:34]
  wire  cout_1367 = cout_1262 & cout_1263; // @[Mul.scala 207:34]
  wire  sum_1368 = sum_1266 ^ sum_1267; // @[Mul.scala 206:34]
  wire  cout_1368 = sum_1266 & sum_1267; // @[Mul.scala 207:34]
  wire  sum_1369 = cout_1264 ^ cout_1265; // @[Mul.scala 206:34]
  wire  cout_1369 = cout_1264 & cout_1265; // @[Mul.scala 207:34]
  wire  sum_1370 = sum_1268 ^ sum_1269; // @[Mul.scala 206:34]
  wire  cout_1370 = sum_1268 & sum_1269; // @[Mul.scala 207:34]
  wire  sum_1371 = cout_1266 ^ cout_1267; // @[Mul.scala 206:34]
  wire  cout_1371 = cout_1266 & cout_1267; // @[Mul.scala 207:34]
  wire  sum_1372 = sum_1270 ^ sum_1271; // @[Mul.scala 206:34]
  wire  cout_1372 = sum_1270 & sum_1271; // @[Mul.scala 207:34]
  wire  sum_1373 = cout_1268 ^ cout_1269; // @[Mul.scala 206:34]
  wire  cout_1373 = cout_1268 & cout_1269; // @[Mul.scala 207:34]
  wire  _sum_T_2000 = sum_1272 ^ cout_1270; // @[Mul.scala 191:34]
  wire  sum_1374 = sum_1272 ^ cout_1270 ^ cout_1271; // @[Mul.scala 191:42]
  wire  cout_1374 = sum_1272 & cout_1270 | _sum_T_2000 & cout_1271; // @[Mul.scala 192:44]
  wire  sum_1375 = sum_1273 ^ cout_1272; // @[Mul.scala 206:34]
  wire  cout_1375 = sum_1273 & cout_1272; // @[Mul.scala 207:34]
  wire  sum_1376 = sum_1274 ^ cout_1273; // @[Mul.scala 206:34]
  wire  cout_1376 = sum_1274 & cout_1273; // @[Mul.scala 207:34]
  wire  sum_1377 = sum_1275 ^ cout_1274; // @[Mul.scala 206:34]
  wire  cout_1377 = sum_1275 & cout_1274; // @[Mul.scala 207:34]
  wire  sum_1378 = sum_1276 ^ cout_1275; // @[Mul.scala 206:34]
  wire  cout_1378 = sum_1276 & cout_1275; // @[Mul.scala 207:34]
  wire  sum_1379 = sum_1277 ^ cout_1276; // @[Mul.scala 206:34]
  wire  sum_1395 = sum_1293 ^ cout_1292; // @[Mul.scala 206:34]
  wire  cout_1395 = sum_1293 & cout_1292; // @[Mul.scala 207:34]
  wire  sum_1396 = sum_1294 ^ cout_1293; // @[Mul.scala 206:34]
  wire  cout_1396 = sum_1294 & cout_1293; // @[Mul.scala 207:34]
  wire  sum_1397 = sum_1295 ^ cout_1294; // @[Mul.scala 206:34]
  wire  cout_1397 = sum_1295 & cout_1294; // @[Mul.scala 207:34]
  wire  _sum_T_2025 = sum_1296 ^ sum_1297; // @[Mul.scala 191:34]
  wire  sum_1398 = sum_1296 ^ sum_1297 ^ cout_1295; // @[Mul.scala 191:42]
  wire  cout_1398 = sum_1296 & sum_1297 | _sum_T_2025 & cout_1295; // @[Mul.scala 192:44]
  wire  sum_1399 = sum_1298 ^ sum_1299; // @[Mul.scala 206:34]
  wire  cout_1399 = sum_1298 & sum_1299; // @[Mul.scala 207:34]
  wire  sum_1400 = cout_1296 ^ cout_1297; // @[Mul.scala 206:34]
  wire  cout_1400 = cout_1296 & cout_1297; // @[Mul.scala 207:34]
  wire  sum_1401 = sum_1300 ^ sum_1301; // @[Mul.scala 206:34]
  wire  cout_1401 = sum_1300 & sum_1301; // @[Mul.scala 207:34]
  wire  sum_1402 = cout_1298 ^ cout_1299; // @[Mul.scala 206:34]
  wire  cout_1402 = cout_1298 & cout_1299; // @[Mul.scala 207:34]
  wire  sum_1403 = sum_1302 ^ sum_1303; // @[Mul.scala 206:34]
  wire  cout_1403 = sum_1302 & sum_1303; // @[Mul.scala 207:34]
  wire  sum_1404 = cout_1300 ^ cout_1301; // @[Mul.scala 206:34]
  wire  cout_1404 = cout_1300 & cout_1301; // @[Mul.scala 207:34]
  wire  sum_1405 = sum_1304 ^ sum_1305; // @[Mul.scala 206:34]
  wire  cout_1405 = sum_1304 & sum_1305; // @[Mul.scala 207:34]
  wire  sum_1406 = cout_1302 ^ cout_1303; // @[Mul.scala 206:34]
  wire  cout_1406 = cout_1302 & cout_1303; // @[Mul.scala 207:34]
  wire  sum_1407 = sum_1306 ^ sum_1307; // @[Mul.scala 206:34]
  wire  cout_1407 = sum_1306 & sum_1307; // @[Mul.scala 207:34]
  wire  sum_1408 = cout_1304 ^ cout_1305; // @[Mul.scala 206:34]
  wire  cout_1408 = cout_1304 & cout_1305; // @[Mul.scala 207:34]
  wire  sum_1409 = sum_1308 ^ sum_1309; // @[Mul.scala 206:34]
  wire  cout_1409 = sum_1308 & sum_1309; // @[Mul.scala 207:34]
  wire  sum_1410 = cout_1306 ^ cout_1307; // @[Mul.scala 206:34]
  wire  cout_1410 = cout_1306 & cout_1307; // @[Mul.scala 207:34]
  wire  sum_1411 = sum_1310 ^ sum_1311; // @[Mul.scala 206:34]
  wire  cout_1411 = sum_1310 & sum_1311; // @[Mul.scala 207:34]
  wire  sum_1412 = cout_1308 ^ cout_1309; // @[Mul.scala 206:34]
  wire  cout_1412 = cout_1308 & cout_1309; // @[Mul.scala 207:34]
  wire  sum_1413 = sum_1312 ^ sum_1313; // @[Mul.scala 206:34]
  wire  cout_1413 = sum_1312 & sum_1313; // @[Mul.scala 207:34]
  wire  sum_1414 = cout_1310 ^ cout_1311; // @[Mul.scala 206:34]
  wire  cout_1414 = cout_1310 & cout_1311; // @[Mul.scala 207:34]
  wire  sum_1415 = sum_1314 ^ sum_1315; // @[Mul.scala 206:34]
  wire  cout_1415 = sum_1314 & sum_1315; // @[Mul.scala 207:34]
  wire  sum_1416 = cout_1312 ^ cout_1313; // @[Mul.scala 206:34]
  wire  cout_1416 = cout_1312 & cout_1313; // @[Mul.scala 207:34]
  wire  sum_1417 = sum_1316 ^ sum_1317; // @[Mul.scala 206:34]
  wire  cout_1417 = sum_1316 & sum_1317; // @[Mul.scala 207:34]
  wire  sum_1418 = cout_1314 ^ cout_1315; // @[Mul.scala 206:34]
  wire  cout_1418 = cout_1314 & cout_1315; // @[Mul.scala 207:34]
  wire  sum_1419 = sum_1318 ^ sum_1319; // @[Mul.scala 206:34]
  wire  cout_1419 = sum_1318 & sum_1319; // @[Mul.scala 207:34]
  wire  sum_1420 = cout_1316 ^ cout_1317; // @[Mul.scala 206:34]
  wire  cout_1420 = cout_1316 & cout_1317; // @[Mul.scala 207:34]
  wire  sum_1421 = sum_1320 ^ sum_1321; // @[Mul.scala 206:34]
  wire  cout_1421 = sum_1320 & sum_1321; // @[Mul.scala 207:34]
  wire  sum_1422 = cout_1318 ^ cout_1319; // @[Mul.scala 206:34]
  wire  cout_1422 = cout_1318 & cout_1319; // @[Mul.scala 207:34]
  wire  sum_1423 = sum_1322 ^ sum_1323; // @[Mul.scala 206:34]
  wire  cout_1423 = sum_1322 & sum_1323; // @[Mul.scala 207:34]
  wire  sum_1424 = cout_1320 ^ cout_1321; // @[Mul.scala 206:34]
  wire  cout_1424 = cout_1320 & cout_1321; // @[Mul.scala 207:34]
  wire  sum_1425 = sum_1324 ^ sum_1325; // @[Mul.scala 206:34]
  wire  cout_1425 = sum_1324 & sum_1325; // @[Mul.scala 207:34]
  wire  sum_1426 = cout_1322 ^ cout_1323; // @[Mul.scala 206:34]
  wire  cout_1426 = cout_1322 & cout_1323; // @[Mul.scala 207:34]
  wire  sum_1427 = sum_1326 ^ sum_1327; // @[Mul.scala 206:34]
  wire  cout_1427 = sum_1326 & sum_1327; // @[Mul.scala 207:34]
  wire  sum_1428 = cout_1324 ^ cout_1325; // @[Mul.scala 206:34]
  wire  cout_1428 = cout_1324 & cout_1325; // @[Mul.scala 207:34]
  wire  sum_1429 = sum_1328 ^ sum_1329; // @[Mul.scala 206:34]
  wire  cout_1429 = sum_1328 & sum_1329; // @[Mul.scala 207:34]
  wire  sum_1430 = cout_1326 ^ cout_1327; // @[Mul.scala 206:34]
  wire  cout_1430 = cout_1326 & cout_1327; // @[Mul.scala 207:34]
  wire  sum_1431 = sum_1330 ^ sum_1331; // @[Mul.scala 206:34]
  wire  cout_1431 = sum_1330 & sum_1331; // @[Mul.scala 207:34]
  wire  sum_1432 = cout_1328 ^ cout_1329; // @[Mul.scala 206:34]
  wire  cout_1432 = cout_1328 & cout_1329; // @[Mul.scala 207:34]
  wire  sum_1433 = sum_1332 ^ sum_1333; // @[Mul.scala 206:34]
  wire  cout_1433 = sum_1332 & sum_1333; // @[Mul.scala 207:34]
  wire  sum_1434 = cout_1330 ^ cout_1331; // @[Mul.scala 206:34]
  wire  cout_1434 = cout_1330 & cout_1331; // @[Mul.scala 207:34]
  wire  sum_1435 = sum_1334 ^ sum_1335; // @[Mul.scala 206:34]
  wire  cout_1435 = sum_1334 & sum_1335; // @[Mul.scala 207:34]
  wire  sum_1436 = cout_1332 ^ cout_1333; // @[Mul.scala 206:34]
  wire  cout_1436 = cout_1332 & cout_1333; // @[Mul.scala 207:34]
  wire  sum_1437 = sum_1336 ^ sum_1337; // @[Mul.scala 206:34]
  wire  cout_1437 = sum_1336 & sum_1337; // @[Mul.scala 207:34]
  wire  sum_1438 = cout_1334 ^ cout_1335; // @[Mul.scala 206:34]
  wire  cout_1438 = cout_1334 & cout_1335; // @[Mul.scala 207:34]
  wire  sum_1439 = sum_1338 ^ sum_1339; // @[Mul.scala 206:34]
  wire  cout_1439 = sum_1338 & sum_1339; // @[Mul.scala 207:34]
  wire  sum_1440 = cout_1336 ^ cout_1337; // @[Mul.scala 206:34]
  wire  cout_1440 = cout_1336 & cout_1337; // @[Mul.scala 207:34]
  wire  sum_1441 = sum_1340 ^ sum_1341; // @[Mul.scala 206:34]
  wire  cout_1441 = sum_1340 & sum_1341; // @[Mul.scala 207:34]
  wire  sum_1442 = cout_1338 ^ cout_1339; // @[Mul.scala 206:34]
  wire  cout_1442 = cout_1338 & cout_1339; // @[Mul.scala 207:34]
  wire  sum_1443 = sum_1342 ^ sum_1343; // @[Mul.scala 206:34]
  wire  cout_1443 = sum_1342 & sum_1343; // @[Mul.scala 207:34]
  wire  sum_1444 = cout_1340 ^ cout_1341; // @[Mul.scala 206:34]
  wire  cout_1444 = cout_1340 & cout_1341; // @[Mul.scala 207:34]
  wire  sum_1445 = sum_1344 ^ sum_1345; // @[Mul.scala 206:34]
  wire  cout_1445 = sum_1344 & sum_1345; // @[Mul.scala 207:34]
  wire  sum_1446 = cout_1342 ^ cout_1343; // @[Mul.scala 206:34]
  wire  cout_1446 = cout_1342 & cout_1343; // @[Mul.scala 207:34]
  wire  sum_1447 = sum_1346 ^ sum_1347; // @[Mul.scala 206:34]
  wire  cout_1447 = sum_1346 & sum_1347; // @[Mul.scala 207:34]
  wire  sum_1448 = cout_1344 ^ cout_1345; // @[Mul.scala 206:34]
  wire  cout_1448 = cout_1344 & cout_1345; // @[Mul.scala 207:34]
  wire  sum_1449 = sum_1348 ^ sum_1349; // @[Mul.scala 206:34]
  wire  cout_1449 = sum_1348 & sum_1349; // @[Mul.scala 207:34]
  wire  sum_1450 = cout_1346 ^ cout_1347; // @[Mul.scala 206:34]
  wire  cout_1450 = cout_1346 & cout_1347; // @[Mul.scala 207:34]
  wire  sum_1451 = sum_1350 ^ sum_1351; // @[Mul.scala 206:34]
  wire  cout_1451 = sum_1350 & sum_1351; // @[Mul.scala 207:34]
  wire  sum_1452 = cout_1348 ^ cout_1349; // @[Mul.scala 206:34]
  wire  cout_1452 = cout_1348 & cout_1349; // @[Mul.scala 207:34]
  wire  sum_1453 = sum_1352 ^ sum_1353; // @[Mul.scala 206:34]
  wire  cout_1453 = sum_1352 & sum_1353; // @[Mul.scala 207:34]
  wire  sum_1454 = cout_1350 ^ cout_1351; // @[Mul.scala 206:34]
  wire  cout_1454 = cout_1350 & cout_1351; // @[Mul.scala 207:34]
  wire  sum_1455 = sum_1354 ^ sum_1355; // @[Mul.scala 206:34]
  wire  cout_1455 = sum_1354 & sum_1355; // @[Mul.scala 207:34]
  wire  sum_1456 = cout_1352 ^ cout_1353; // @[Mul.scala 206:34]
  wire  cout_1456 = cout_1352 & cout_1353; // @[Mul.scala 207:34]
  wire  sum_1457 = sum_1356 ^ sum_1357; // @[Mul.scala 206:34]
  wire  cout_1457 = sum_1356 & sum_1357; // @[Mul.scala 207:34]
  wire  sum_1458 = cout_1354 ^ cout_1355; // @[Mul.scala 206:34]
  wire  cout_1458 = cout_1354 & cout_1355; // @[Mul.scala 207:34]
  wire  sum_1459 = sum_1358 ^ sum_1359; // @[Mul.scala 206:34]
  wire  cout_1459 = sum_1358 & sum_1359; // @[Mul.scala 207:34]
  wire  sum_1460 = cout_1356 ^ cout_1357; // @[Mul.scala 206:34]
  wire  cout_1460 = cout_1356 & cout_1357; // @[Mul.scala 207:34]
  wire  sum_1461 = sum_1360 ^ sum_1361; // @[Mul.scala 206:34]
  wire  cout_1461 = sum_1360 & sum_1361; // @[Mul.scala 207:34]
  wire  sum_1462 = cout_1358 ^ cout_1359; // @[Mul.scala 206:34]
  wire  cout_1462 = cout_1358 & cout_1359; // @[Mul.scala 207:34]
  wire  sum_1463 = sum_1362 ^ sum_1363; // @[Mul.scala 206:34]
  wire  cout_1463 = sum_1362 & sum_1363; // @[Mul.scala 207:34]
  wire  sum_1464 = cout_1360 ^ cout_1361; // @[Mul.scala 206:34]
  wire  cout_1464 = cout_1360 & cout_1361; // @[Mul.scala 207:34]
  wire  sum_1465 = sum_1364 ^ sum_1365; // @[Mul.scala 206:34]
  wire  cout_1465 = sum_1364 & sum_1365; // @[Mul.scala 207:34]
  wire  sum_1466 = cout_1362 ^ cout_1363; // @[Mul.scala 206:34]
  wire  cout_1466 = cout_1362 & cout_1363; // @[Mul.scala 207:34]
  wire  sum_1467 = sum_1366 ^ sum_1367; // @[Mul.scala 206:34]
  wire  cout_1467 = sum_1366 & sum_1367; // @[Mul.scala 207:34]
  wire  sum_1468 = cout_1364 ^ cout_1365; // @[Mul.scala 206:34]
  wire  cout_1468 = cout_1364 & cout_1365; // @[Mul.scala 207:34]
  wire  sum_1469 = sum_1368 ^ sum_1369; // @[Mul.scala 206:34]
  wire  cout_1469 = sum_1368 & sum_1369; // @[Mul.scala 207:34]
  wire  sum_1470 = cout_1366 ^ cout_1367; // @[Mul.scala 206:34]
  wire  cout_1470 = cout_1366 & cout_1367; // @[Mul.scala 207:34]
  wire  sum_1471 = sum_1370 ^ sum_1371; // @[Mul.scala 206:34]
  wire  cout_1471 = sum_1370 & sum_1371; // @[Mul.scala 207:34]
  wire  sum_1472 = cout_1368 ^ cout_1369; // @[Mul.scala 206:34]
  wire  cout_1472 = cout_1368 & cout_1369; // @[Mul.scala 207:34]
  wire  sum_1473 = sum_1372 ^ sum_1373; // @[Mul.scala 206:34]
  wire  cout_1473 = sum_1372 & sum_1373; // @[Mul.scala 207:34]
  wire  sum_1474 = cout_1370 ^ cout_1371; // @[Mul.scala 206:34]
  wire  cout_1474 = cout_1370 & cout_1371; // @[Mul.scala 207:34]
  wire  _sum_T_2103 = sum_1374 ^ cout_1372; // @[Mul.scala 191:34]
  wire  sum_1475 = sum_1374 ^ cout_1372 ^ cout_1373; // @[Mul.scala 191:42]
  wire  cout_1475 = sum_1374 & cout_1372 | _sum_T_2103 & cout_1373; // @[Mul.scala 192:44]
  wire  sum_1476 = sum_1375 ^ cout_1374; // @[Mul.scala 206:34]
  wire  cout_1476 = sum_1375 & cout_1374; // @[Mul.scala 207:34]
  wire  sum_1477 = sum_1376 ^ cout_1375; // @[Mul.scala 206:34]
  wire  cout_1477 = sum_1376 & cout_1375; // @[Mul.scala 207:34]
  wire  sum_1478 = sum_1377 ^ cout_1376; // @[Mul.scala 206:34]
  wire  cout_1478 = sum_1377 & cout_1376; // @[Mul.scala 207:34]
  wire  sum_1479 = sum_1378 ^ cout_1377; // @[Mul.scala 206:34]
  wire  cout_1479 = sum_1378 & cout_1377; // @[Mul.scala 207:34]
  wire  sum_1480 = sum_1379 ^ cout_1378; // @[Mul.scala 206:34]
  wire  sum_1497 = sum_1396 ^ cout_1395; // @[Mul.scala 206:34]
  wire  cout_1497 = sum_1396 & cout_1395; // @[Mul.scala 207:34]
  wire  sum_1498 = sum_1397 ^ cout_1396; // @[Mul.scala 206:34]
  wire  cout_1498 = sum_1397 & cout_1396; // @[Mul.scala 207:34]
  wire  sum_1499 = sum_1398 ^ cout_1397; // @[Mul.scala 206:34]
  wire  cout_1499 = sum_1398 & cout_1397; // @[Mul.scala 207:34]
  wire  _sum_T_2129 = sum_1399 ^ sum_1400; // @[Mul.scala 191:34]
  wire  sum_1500 = sum_1399 ^ sum_1400 ^ cout_1398; // @[Mul.scala 191:42]
  wire  cout_1500 = sum_1399 & sum_1400 | _sum_T_2129 & cout_1398; // @[Mul.scala 192:44]
  wire  sum_1501 = sum_1401 ^ sum_1402; // @[Mul.scala 206:34]
  wire  cout_1501 = sum_1401 & sum_1402; // @[Mul.scala 207:34]
  wire  sum_1502 = cout_1399 ^ cout_1400; // @[Mul.scala 206:34]
  wire  cout_1502 = cout_1399 & cout_1400; // @[Mul.scala 207:34]
  wire  sum_1503 = sum_1403 ^ sum_1404; // @[Mul.scala 206:34]
  wire  cout_1503 = sum_1403 & sum_1404; // @[Mul.scala 207:34]
  wire  sum_1504 = cout_1401 ^ cout_1402; // @[Mul.scala 206:34]
  wire  cout_1504 = cout_1401 & cout_1402; // @[Mul.scala 207:34]
  wire  sum_1505 = sum_1405 ^ sum_1406; // @[Mul.scala 206:34]
  wire  cout_1505 = sum_1405 & sum_1406; // @[Mul.scala 207:34]
  wire  sum_1506 = cout_1403 ^ cout_1404; // @[Mul.scala 206:34]
  wire  cout_1506 = cout_1403 & cout_1404; // @[Mul.scala 207:34]
  wire  sum_1507 = sum_1407 ^ sum_1408; // @[Mul.scala 206:34]
  wire  cout_1507 = sum_1407 & sum_1408; // @[Mul.scala 207:34]
  wire  sum_1508 = cout_1405 ^ cout_1406; // @[Mul.scala 206:34]
  wire  cout_1508 = cout_1405 & cout_1406; // @[Mul.scala 207:34]
  wire  sum_1509 = sum_1409 ^ sum_1410; // @[Mul.scala 206:34]
  wire  cout_1509 = sum_1409 & sum_1410; // @[Mul.scala 207:34]
  wire  sum_1510 = cout_1407 ^ cout_1408; // @[Mul.scala 206:34]
  wire  cout_1510 = cout_1407 & cout_1408; // @[Mul.scala 207:34]
  wire  sum_1511 = sum_1411 ^ sum_1412; // @[Mul.scala 206:34]
  wire  cout_1511 = sum_1411 & sum_1412; // @[Mul.scala 207:34]
  wire  sum_1512 = cout_1409 ^ cout_1410; // @[Mul.scala 206:34]
  wire  cout_1512 = cout_1409 & cout_1410; // @[Mul.scala 207:34]
  wire  sum_1513 = sum_1413 ^ sum_1414; // @[Mul.scala 206:34]
  wire  cout_1513 = sum_1413 & sum_1414; // @[Mul.scala 207:34]
  wire  sum_1514 = cout_1411 ^ cout_1412; // @[Mul.scala 206:34]
  wire  cout_1514 = cout_1411 & cout_1412; // @[Mul.scala 207:34]
  wire  sum_1515 = sum_1415 ^ sum_1416; // @[Mul.scala 206:34]
  wire  cout_1515 = sum_1415 & sum_1416; // @[Mul.scala 207:34]
  wire  sum_1516 = cout_1413 ^ cout_1414; // @[Mul.scala 206:34]
  wire  cout_1516 = cout_1413 & cout_1414; // @[Mul.scala 207:34]
  wire  sum_1517 = sum_1417 ^ sum_1418; // @[Mul.scala 206:34]
  wire  cout_1517 = sum_1417 & sum_1418; // @[Mul.scala 207:34]
  wire  sum_1518 = cout_1415 ^ cout_1416; // @[Mul.scala 206:34]
  wire  cout_1518 = cout_1415 & cout_1416; // @[Mul.scala 207:34]
  wire  sum_1519 = sum_1419 ^ sum_1420; // @[Mul.scala 206:34]
  wire  cout_1519 = sum_1419 & sum_1420; // @[Mul.scala 207:34]
  wire  sum_1520 = cout_1417 ^ cout_1418; // @[Mul.scala 206:34]
  wire  cout_1520 = cout_1417 & cout_1418; // @[Mul.scala 207:34]
  wire  sum_1521 = sum_1421 ^ sum_1422; // @[Mul.scala 206:34]
  wire  cout_1521 = sum_1421 & sum_1422; // @[Mul.scala 207:34]
  wire  sum_1522 = cout_1419 ^ cout_1420; // @[Mul.scala 206:34]
  wire  cout_1522 = cout_1419 & cout_1420; // @[Mul.scala 207:34]
  wire  sum_1523 = sum_1423 ^ sum_1424; // @[Mul.scala 206:34]
  wire  cout_1523 = sum_1423 & sum_1424; // @[Mul.scala 207:34]
  wire  sum_1524 = cout_1421 ^ cout_1422; // @[Mul.scala 206:34]
  wire  cout_1524 = cout_1421 & cout_1422; // @[Mul.scala 207:34]
  wire  sum_1525 = sum_1425 ^ sum_1426; // @[Mul.scala 206:34]
  wire  cout_1525 = sum_1425 & sum_1426; // @[Mul.scala 207:34]
  wire  sum_1526 = cout_1423 ^ cout_1424; // @[Mul.scala 206:34]
  wire  cout_1526 = cout_1423 & cout_1424; // @[Mul.scala 207:34]
  wire  sum_1527 = sum_1427 ^ sum_1428; // @[Mul.scala 206:34]
  wire  cout_1527 = sum_1427 & sum_1428; // @[Mul.scala 207:34]
  wire  sum_1528 = cout_1425 ^ cout_1426; // @[Mul.scala 206:34]
  wire  cout_1528 = cout_1425 & cout_1426; // @[Mul.scala 207:34]
  wire  sum_1529 = sum_1429 ^ sum_1430; // @[Mul.scala 206:34]
  wire  cout_1529 = sum_1429 & sum_1430; // @[Mul.scala 207:34]
  wire  sum_1530 = cout_1427 ^ cout_1428; // @[Mul.scala 206:34]
  wire  cout_1530 = cout_1427 & cout_1428; // @[Mul.scala 207:34]
  wire  sum_1531 = sum_1431 ^ sum_1432; // @[Mul.scala 206:34]
  wire  cout_1531 = sum_1431 & sum_1432; // @[Mul.scala 207:34]
  wire  sum_1532 = cout_1429 ^ cout_1430; // @[Mul.scala 206:34]
  wire  cout_1532 = cout_1429 & cout_1430; // @[Mul.scala 207:34]
  wire  sum_1533 = sum_1433 ^ sum_1434; // @[Mul.scala 206:34]
  wire  cout_1533 = sum_1433 & sum_1434; // @[Mul.scala 207:34]
  wire  sum_1534 = cout_1431 ^ cout_1432; // @[Mul.scala 206:34]
  wire  cout_1534 = cout_1431 & cout_1432; // @[Mul.scala 207:34]
  wire  sum_1535 = sum_1435 ^ sum_1436; // @[Mul.scala 206:34]
  wire  cout_1535 = sum_1435 & sum_1436; // @[Mul.scala 207:34]
  wire  sum_1536 = cout_1433 ^ cout_1434; // @[Mul.scala 206:34]
  wire  cout_1536 = cout_1433 & cout_1434; // @[Mul.scala 207:34]
  wire  sum_1537 = sum_1437 ^ sum_1438; // @[Mul.scala 206:34]
  wire  cout_1537 = sum_1437 & sum_1438; // @[Mul.scala 207:34]
  wire  sum_1538 = cout_1435 ^ cout_1436; // @[Mul.scala 206:34]
  wire  cout_1538 = cout_1435 & cout_1436; // @[Mul.scala 207:34]
  wire  sum_1539 = sum_1439 ^ sum_1440; // @[Mul.scala 206:34]
  wire  cout_1539 = sum_1439 & sum_1440; // @[Mul.scala 207:34]
  wire  sum_1540 = cout_1437 ^ cout_1438; // @[Mul.scala 206:34]
  wire  cout_1540 = cout_1437 & cout_1438; // @[Mul.scala 207:34]
  wire  sum_1541 = sum_1441 ^ sum_1442; // @[Mul.scala 206:34]
  wire  cout_1541 = sum_1441 & sum_1442; // @[Mul.scala 207:34]
  wire  sum_1542 = cout_1439 ^ cout_1440; // @[Mul.scala 206:34]
  wire  cout_1542 = cout_1439 & cout_1440; // @[Mul.scala 207:34]
  wire  sum_1543 = sum_1443 ^ sum_1444; // @[Mul.scala 206:34]
  wire  cout_1543 = sum_1443 & sum_1444; // @[Mul.scala 207:34]
  wire  sum_1544 = cout_1441 ^ cout_1442; // @[Mul.scala 206:34]
  wire  cout_1544 = cout_1441 & cout_1442; // @[Mul.scala 207:34]
  wire  sum_1545 = sum_1445 ^ sum_1446; // @[Mul.scala 206:34]
  wire  cout_1545 = sum_1445 & sum_1446; // @[Mul.scala 207:34]
  wire  sum_1546 = cout_1443 ^ cout_1444; // @[Mul.scala 206:34]
  wire  cout_1546 = cout_1443 & cout_1444; // @[Mul.scala 207:34]
  wire  sum_1547 = sum_1447 ^ sum_1448; // @[Mul.scala 206:34]
  wire  cout_1547 = sum_1447 & sum_1448; // @[Mul.scala 207:34]
  wire  sum_1548 = cout_1445 ^ cout_1446; // @[Mul.scala 206:34]
  wire  cout_1548 = cout_1445 & cout_1446; // @[Mul.scala 207:34]
  wire  sum_1549 = sum_1449 ^ sum_1450; // @[Mul.scala 206:34]
  wire  cout_1549 = sum_1449 & sum_1450; // @[Mul.scala 207:34]
  wire  sum_1550 = cout_1447 ^ cout_1448; // @[Mul.scala 206:34]
  wire  cout_1550 = cout_1447 & cout_1448; // @[Mul.scala 207:34]
  wire  sum_1551 = sum_1451 ^ sum_1452; // @[Mul.scala 206:34]
  wire  cout_1551 = sum_1451 & sum_1452; // @[Mul.scala 207:34]
  wire  sum_1552 = cout_1449 ^ cout_1450; // @[Mul.scala 206:34]
  wire  cout_1552 = cout_1449 & cout_1450; // @[Mul.scala 207:34]
  wire  sum_1553 = sum_1453 ^ sum_1454; // @[Mul.scala 206:34]
  wire  cout_1553 = sum_1453 & sum_1454; // @[Mul.scala 207:34]
  wire  sum_1554 = cout_1451 ^ cout_1452; // @[Mul.scala 206:34]
  wire  cout_1554 = cout_1451 & cout_1452; // @[Mul.scala 207:34]
  wire  sum_1555 = sum_1455 ^ sum_1456; // @[Mul.scala 206:34]
  wire  cout_1555 = sum_1455 & sum_1456; // @[Mul.scala 207:34]
  wire  sum_1556 = cout_1453 ^ cout_1454; // @[Mul.scala 206:34]
  wire  cout_1556 = cout_1453 & cout_1454; // @[Mul.scala 207:34]
  wire  sum_1557 = sum_1457 ^ sum_1458; // @[Mul.scala 206:34]
  wire  cout_1557 = sum_1457 & sum_1458; // @[Mul.scala 207:34]
  wire  sum_1558 = cout_1455 ^ cout_1456; // @[Mul.scala 206:34]
  wire  cout_1558 = cout_1455 & cout_1456; // @[Mul.scala 207:34]
  wire  sum_1559 = sum_1459 ^ sum_1460; // @[Mul.scala 206:34]
  wire  cout_1559 = sum_1459 & sum_1460; // @[Mul.scala 207:34]
  wire  sum_1560 = cout_1457 ^ cout_1458; // @[Mul.scala 206:34]
  wire  cout_1560 = cout_1457 & cout_1458; // @[Mul.scala 207:34]
  wire  sum_1561 = sum_1461 ^ sum_1462; // @[Mul.scala 206:34]
  wire  cout_1561 = sum_1461 & sum_1462; // @[Mul.scala 207:34]
  wire  sum_1562 = cout_1459 ^ cout_1460; // @[Mul.scala 206:34]
  wire  cout_1562 = cout_1459 & cout_1460; // @[Mul.scala 207:34]
  wire  sum_1563 = sum_1463 ^ sum_1464; // @[Mul.scala 206:34]
  wire  cout_1563 = sum_1463 & sum_1464; // @[Mul.scala 207:34]
  wire  sum_1564 = cout_1461 ^ cout_1462; // @[Mul.scala 206:34]
  wire  cout_1564 = cout_1461 & cout_1462; // @[Mul.scala 207:34]
  wire  sum_1565 = sum_1465 ^ sum_1466; // @[Mul.scala 206:34]
  wire  cout_1565 = sum_1465 & sum_1466; // @[Mul.scala 207:34]
  wire  sum_1566 = cout_1463 ^ cout_1464; // @[Mul.scala 206:34]
  wire  cout_1566 = cout_1463 & cout_1464; // @[Mul.scala 207:34]
  wire  sum_1567 = sum_1467 ^ sum_1468; // @[Mul.scala 206:34]
  wire  cout_1567 = sum_1467 & sum_1468; // @[Mul.scala 207:34]
  wire  sum_1568 = cout_1465 ^ cout_1466; // @[Mul.scala 206:34]
  wire  cout_1568 = cout_1465 & cout_1466; // @[Mul.scala 207:34]
  wire  sum_1569 = sum_1469 ^ sum_1470; // @[Mul.scala 206:34]
  wire  cout_1569 = sum_1469 & sum_1470; // @[Mul.scala 207:34]
  wire  sum_1570 = cout_1467 ^ cout_1468; // @[Mul.scala 206:34]
  wire  cout_1570 = cout_1467 & cout_1468; // @[Mul.scala 207:34]
  wire  sum_1571 = sum_1471 ^ sum_1472; // @[Mul.scala 206:34]
  wire  cout_1571 = sum_1471 & sum_1472; // @[Mul.scala 207:34]
  wire  sum_1572 = cout_1469 ^ cout_1470; // @[Mul.scala 206:34]
  wire  cout_1572 = cout_1469 & cout_1470; // @[Mul.scala 207:34]
  wire  sum_1573 = sum_1473 ^ sum_1474; // @[Mul.scala 206:34]
  wire  cout_1573 = sum_1473 & sum_1474; // @[Mul.scala 207:34]
  wire  sum_1574 = cout_1471 ^ cout_1472; // @[Mul.scala 206:34]
  wire  cout_1574 = cout_1471 & cout_1472; // @[Mul.scala 207:34]
  wire  _sum_T_2205 = sum_1475 ^ cout_1473; // @[Mul.scala 191:34]
  wire  sum_1575 = sum_1475 ^ cout_1473 ^ cout_1474; // @[Mul.scala 191:42]
  wire  cout_1575 = sum_1475 & cout_1473 | _sum_T_2205 & cout_1474; // @[Mul.scala 192:44]
  wire  sum_1576 = sum_1476 ^ cout_1475; // @[Mul.scala 206:34]
  wire  cout_1576 = sum_1476 & cout_1475; // @[Mul.scala 207:34]
  wire  sum_1577 = sum_1477 ^ cout_1476; // @[Mul.scala 206:34]
  wire  cout_1577 = sum_1477 & cout_1476; // @[Mul.scala 207:34]
  wire  sum_1578 = sum_1478 ^ cout_1477; // @[Mul.scala 206:34]
  wire  cout_1578 = sum_1478 & cout_1477; // @[Mul.scala 207:34]
  wire  sum_1579 = sum_1479 ^ cout_1478; // @[Mul.scala 206:34]
  wire  cout_1579 = sum_1479 & cout_1478; // @[Mul.scala 207:34]
  wire  sum_1580 = sum_1480 ^ cout_1479; // @[Mul.scala 206:34]
  wire  sum_1598 = sum_1498 ^ cout_1497; // @[Mul.scala 206:34]
  wire  cout_1598 = sum_1498 & cout_1497; // @[Mul.scala 207:34]
  wire  sum_1599 = sum_1499 ^ cout_1498; // @[Mul.scala 206:34]
  wire  cout_1599 = sum_1499 & cout_1498; // @[Mul.scala 207:34]
  wire  sum_1600 = sum_1500 ^ cout_1499; // @[Mul.scala 206:34]
  wire  cout_1600 = sum_1500 & cout_1499; // @[Mul.scala 207:34]
  wire  _sum_T_2232 = sum_1501 ^ sum_1502; // @[Mul.scala 191:34]
  wire  sum_1601 = sum_1501 ^ sum_1502 ^ cout_1500; // @[Mul.scala 191:42]
  wire  cout_1601 = sum_1501 & sum_1502 | _sum_T_2232 & cout_1500; // @[Mul.scala 192:44]
  wire  sum_1602 = sum_1503 ^ sum_1504; // @[Mul.scala 206:34]
  wire  cout_1602 = sum_1503 & sum_1504; // @[Mul.scala 207:34]
  wire  sum_1603 = cout_1501 ^ cout_1502; // @[Mul.scala 206:34]
  wire  cout_1603 = cout_1501 & cout_1502; // @[Mul.scala 207:34]
  wire  sum_1604 = sum_1505 ^ sum_1506; // @[Mul.scala 206:34]
  wire  cout_1604 = sum_1505 & sum_1506; // @[Mul.scala 207:34]
  wire  sum_1605 = cout_1503 ^ cout_1504; // @[Mul.scala 206:34]
  wire  cout_1605 = cout_1503 & cout_1504; // @[Mul.scala 207:34]
  wire  sum_1606 = sum_1507 ^ sum_1508; // @[Mul.scala 206:34]
  wire  cout_1606 = sum_1507 & sum_1508; // @[Mul.scala 207:34]
  wire  sum_1607 = cout_1505 ^ cout_1506; // @[Mul.scala 206:34]
  wire  cout_1607 = cout_1505 & cout_1506; // @[Mul.scala 207:34]
  wire  sum_1608 = sum_1509 ^ sum_1510; // @[Mul.scala 206:34]
  wire  cout_1608 = sum_1509 & sum_1510; // @[Mul.scala 207:34]
  wire  sum_1609 = cout_1507 ^ cout_1508; // @[Mul.scala 206:34]
  wire  cout_1609 = cout_1507 & cout_1508; // @[Mul.scala 207:34]
  wire  sum_1610 = sum_1511 ^ sum_1512; // @[Mul.scala 206:34]
  wire  cout_1610 = sum_1511 & sum_1512; // @[Mul.scala 207:34]
  wire  sum_1611 = cout_1509 ^ cout_1510; // @[Mul.scala 206:34]
  wire  cout_1611 = cout_1509 & cout_1510; // @[Mul.scala 207:34]
  wire  sum_1612 = sum_1513 ^ sum_1514; // @[Mul.scala 206:34]
  wire  cout_1612 = sum_1513 & sum_1514; // @[Mul.scala 207:34]
  wire  sum_1613 = cout_1511 ^ cout_1512; // @[Mul.scala 206:34]
  wire  cout_1613 = cout_1511 & cout_1512; // @[Mul.scala 207:34]
  wire  sum_1614 = sum_1515 ^ sum_1516; // @[Mul.scala 206:34]
  wire  cout_1614 = sum_1515 & sum_1516; // @[Mul.scala 207:34]
  wire  sum_1615 = cout_1513 ^ cout_1514; // @[Mul.scala 206:34]
  wire  cout_1615 = cout_1513 & cout_1514; // @[Mul.scala 207:34]
  wire  sum_1616 = sum_1517 ^ sum_1518; // @[Mul.scala 206:34]
  wire  cout_1616 = sum_1517 & sum_1518; // @[Mul.scala 207:34]
  wire  sum_1617 = cout_1515 ^ cout_1516; // @[Mul.scala 206:34]
  wire  cout_1617 = cout_1515 & cout_1516; // @[Mul.scala 207:34]
  wire  sum_1618 = sum_1519 ^ sum_1520; // @[Mul.scala 206:34]
  wire  cout_1618 = sum_1519 & sum_1520; // @[Mul.scala 207:34]
  wire  sum_1619 = cout_1517 ^ cout_1518; // @[Mul.scala 206:34]
  wire  cout_1619 = cout_1517 & cout_1518; // @[Mul.scala 207:34]
  wire  sum_1620 = sum_1521 ^ sum_1522; // @[Mul.scala 206:34]
  wire  cout_1620 = sum_1521 & sum_1522; // @[Mul.scala 207:34]
  wire  sum_1621 = cout_1519 ^ cout_1520; // @[Mul.scala 206:34]
  wire  cout_1621 = cout_1519 & cout_1520; // @[Mul.scala 207:34]
  wire  sum_1622 = sum_1523 ^ sum_1524; // @[Mul.scala 206:34]
  wire  cout_1622 = sum_1523 & sum_1524; // @[Mul.scala 207:34]
  wire  sum_1623 = cout_1521 ^ cout_1522; // @[Mul.scala 206:34]
  wire  cout_1623 = cout_1521 & cout_1522; // @[Mul.scala 207:34]
  wire  sum_1624 = sum_1525 ^ sum_1526; // @[Mul.scala 206:34]
  wire  cout_1624 = sum_1525 & sum_1526; // @[Mul.scala 207:34]
  wire  sum_1625 = cout_1523 ^ cout_1524; // @[Mul.scala 206:34]
  wire  cout_1625 = cout_1523 & cout_1524; // @[Mul.scala 207:34]
  wire  sum_1626 = sum_1527 ^ sum_1528; // @[Mul.scala 206:34]
  wire  cout_1626 = sum_1527 & sum_1528; // @[Mul.scala 207:34]
  wire  sum_1627 = cout_1525 ^ cout_1526; // @[Mul.scala 206:34]
  wire  cout_1627 = cout_1525 & cout_1526; // @[Mul.scala 207:34]
  wire  sum_1628 = sum_1529 ^ sum_1530; // @[Mul.scala 206:34]
  wire  cout_1628 = sum_1529 & sum_1530; // @[Mul.scala 207:34]
  wire  sum_1629 = cout_1527 ^ cout_1528; // @[Mul.scala 206:34]
  wire  cout_1629 = cout_1527 & cout_1528; // @[Mul.scala 207:34]
  wire  sum_1630 = sum_1531 ^ sum_1532; // @[Mul.scala 206:34]
  wire  cout_1630 = sum_1531 & sum_1532; // @[Mul.scala 207:34]
  wire  sum_1631 = cout_1529 ^ cout_1530; // @[Mul.scala 206:34]
  wire  cout_1631 = cout_1529 & cout_1530; // @[Mul.scala 207:34]
  wire  sum_1632 = sum_1533 ^ sum_1534; // @[Mul.scala 206:34]
  wire  cout_1632 = sum_1533 & sum_1534; // @[Mul.scala 207:34]
  wire  sum_1633 = cout_1531 ^ cout_1532; // @[Mul.scala 206:34]
  wire  cout_1633 = cout_1531 & cout_1532; // @[Mul.scala 207:34]
  wire  sum_1634 = sum_1535 ^ sum_1536; // @[Mul.scala 206:34]
  wire  cout_1634 = sum_1535 & sum_1536; // @[Mul.scala 207:34]
  wire  sum_1635 = cout_1533 ^ cout_1534; // @[Mul.scala 206:34]
  wire  cout_1635 = cout_1533 & cout_1534; // @[Mul.scala 207:34]
  wire  sum_1636 = sum_1537 ^ sum_1538; // @[Mul.scala 206:34]
  wire  cout_1636 = sum_1537 & sum_1538; // @[Mul.scala 207:34]
  wire  sum_1637 = cout_1535 ^ cout_1536; // @[Mul.scala 206:34]
  wire  cout_1637 = cout_1535 & cout_1536; // @[Mul.scala 207:34]
  wire  sum_1638 = sum_1539 ^ sum_1540; // @[Mul.scala 206:34]
  wire  cout_1638 = sum_1539 & sum_1540; // @[Mul.scala 207:34]
  wire  sum_1639 = cout_1537 ^ cout_1538; // @[Mul.scala 206:34]
  wire  cout_1639 = cout_1537 & cout_1538; // @[Mul.scala 207:34]
  wire  sum_1640 = sum_1541 ^ sum_1542; // @[Mul.scala 206:34]
  wire  cout_1640 = sum_1541 & sum_1542; // @[Mul.scala 207:34]
  wire  sum_1641 = cout_1539 ^ cout_1540; // @[Mul.scala 206:34]
  wire  cout_1641 = cout_1539 & cout_1540; // @[Mul.scala 207:34]
  wire  sum_1642 = sum_1543 ^ sum_1544; // @[Mul.scala 206:34]
  wire  cout_1642 = sum_1543 & sum_1544; // @[Mul.scala 207:34]
  wire  sum_1643 = cout_1541 ^ cout_1542; // @[Mul.scala 206:34]
  wire  cout_1643 = cout_1541 & cout_1542; // @[Mul.scala 207:34]
  wire  sum_1644 = sum_1545 ^ sum_1546; // @[Mul.scala 206:34]
  wire  cout_1644 = sum_1545 & sum_1546; // @[Mul.scala 207:34]
  wire  sum_1645 = cout_1543 ^ cout_1544; // @[Mul.scala 206:34]
  wire  cout_1645 = cout_1543 & cout_1544; // @[Mul.scala 207:34]
  wire  sum_1646 = sum_1547 ^ sum_1548; // @[Mul.scala 206:34]
  wire  cout_1646 = sum_1547 & sum_1548; // @[Mul.scala 207:34]
  wire  sum_1647 = cout_1545 ^ cout_1546; // @[Mul.scala 206:34]
  wire  cout_1647 = cout_1545 & cout_1546; // @[Mul.scala 207:34]
  wire  sum_1648 = sum_1549 ^ sum_1550; // @[Mul.scala 206:34]
  wire  cout_1648 = sum_1549 & sum_1550; // @[Mul.scala 207:34]
  wire  sum_1649 = cout_1547 ^ cout_1548; // @[Mul.scala 206:34]
  wire  cout_1649 = cout_1547 & cout_1548; // @[Mul.scala 207:34]
  wire  sum_1650 = sum_1551 ^ sum_1552; // @[Mul.scala 206:34]
  wire  cout_1650 = sum_1551 & sum_1552; // @[Mul.scala 207:34]
  wire  sum_1651 = cout_1549 ^ cout_1550; // @[Mul.scala 206:34]
  wire  cout_1651 = cout_1549 & cout_1550; // @[Mul.scala 207:34]
  wire  sum_1652 = sum_1553 ^ sum_1554; // @[Mul.scala 206:34]
  wire  cout_1652 = sum_1553 & sum_1554; // @[Mul.scala 207:34]
  wire  sum_1653 = cout_1551 ^ cout_1552; // @[Mul.scala 206:34]
  wire  cout_1653 = cout_1551 & cout_1552; // @[Mul.scala 207:34]
  wire  sum_1654 = sum_1555 ^ sum_1556; // @[Mul.scala 206:34]
  wire  cout_1654 = sum_1555 & sum_1556; // @[Mul.scala 207:34]
  wire  sum_1655 = cout_1553 ^ cout_1554; // @[Mul.scala 206:34]
  wire  cout_1655 = cout_1553 & cout_1554; // @[Mul.scala 207:34]
  wire  sum_1656 = sum_1557 ^ sum_1558; // @[Mul.scala 206:34]
  wire  cout_1656 = sum_1557 & sum_1558; // @[Mul.scala 207:34]
  wire  sum_1657 = cout_1555 ^ cout_1556; // @[Mul.scala 206:34]
  wire  cout_1657 = cout_1555 & cout_1556; // @[Mul.scala 207:34]
  wire  sum_1658 = sum_1559 ^ sum_1560; // @[Mul.scala 206:34]
  wire  cout_1658 = sum_1559 & sum_1560; // @[Mul.scala 207:34]
  wire  sum_1659 = cout_1557 ^ cout_1558; // @[Mul.scala 206:34]
  wire  cout_1659 = cout_1557 & cout_1558; // @[Mul.scala 207:34]
  wire  sum_1660 = sum_1561 ^ sum_1562; // @[Mul.scala 206:34]
  wire  cout_1660 = sum_1561 & sum_1562; // @[Mul.scala 207:34]
  wire  sum_1661 = cout_1559 ^ cout_1560; // @[Mul.scala 206:34]
  wire  cout_1661 = cout_1559 & cout_1560; // @[Mul.scala 207:34]
  wire  sum_1662 = sum_1563 ^ sum_1564; // @[Mul.scala 206:34]
  wire  cout_1662 = sum_1563 & sum_1564; // @[Mul.scala 207:34]
  wire  sum_1663 = cout_1561 ^ cout_1562; // @[Mul.scala 206:34]
  wire  cout_1663 = cout_1561 & cout_1562; // @[Mul.scala 207:34]
  wire  sum_1664 = sum_1565 ^ sum_1566; // @[Mul.scala 206:34]
  wire  cout_1664 = sum_1565 & sum_1566; // @[Mul.scala 207:34]
  wire  sum_1665 = cout_1563 ^ cout_1564; // @[Mul.scala 206:34]
  wire  cout_1665 = cout_1563 & cout_1564; // @[Mul.scala 207:34]
  wire  sum_1666 = sum_1567 ^ sum_1568; // @[Mul.scala 206:34]
  wire  cout_1666 = sum_1567 & sum_1568; // @[Mul.scala 207:34]
  wire  sum_1667 = cout_1565 ^ cout_1566; // @[Mul.scala 206:34]
  wire  cout_1667 = cout_1565 & cout_1566; // @[Mul.scala 207:34]
  wire  sum_1668 = sum_1569 ^ sum_1570; // @[Mul.scala 206:34]
  wire  cout_1668 = sum_1569 & sum_1570; // @[Mul.scala 207:34]
  wire  sum_1669 = cout_1567 ^ cout_1568; // @[Mul.scala 206:34]
  wire  cout_1669 = cout_1567 & cout_1568; // @[Mul.scala 207:34]
  wire  sum_1670 = sum_1571 ^ sum_1572; // @[Mul.scala 206:34]
  wire  cout_1670 = sum_1571 & sum_1572; // @[Mul.scala 207:34]
  wire  sum_1671 = cout_1569 ^ cout_1570; // @[Mul.scala 206:34]
  wire  cout_1671 = cout_1569 & cout_1570; // @[Mul.scala 207:34]
  wire  sum_1672 = sum_1573 ^ sum_1574; // @[Mul.scala 206:34]
  wire  cout_1672 = sum_1573 & sum_1574; // @[Mul.scala 207:34]
  wire  sum_1673 = cout_1571 ^ cout_1572; // @[Mul.scala 206:34]
  wire  cout_1673 = cout_1571 & cout_1572; // @[Mul.scala 207:34]
  wire  _sum_T_2306 = sum_1575 ^ cout_1573; // @[Mul.scala 191:34]
  wire  sum_1674 = sum_1575 ^ cout_1573 ^ cout_1574; // @[Mul.scala 191:42]
  wire  cout_1674 = sum_1575 & cout_1573 | _sum_T_2306 & cout_1574; // @[Mul.scala 192:44]
  wire  sum_1675 = sum_1576 ^ cout_1575; // @[Mul.scala 206:34]
  wire  cout_1675 = sum_1576 & cout_1575; // @[Mul.scala 207:34]
  wire  sum_1676 = sum_1577 ^ cout_1576; // @[Mul.scala 206:34]
  wire  cout_1676 = sum_1577 & cout_1576; // @[Mul.scala 207:34]
  wire  sum_1677 = sum_1578 ^ cout_1577; // @[Mul.scala 206:34]
  wire  cout_1677 = sum_1578 & cout_1577; // @[Mul.scala 207:34]
  wire  sum_1678 = sum_1579 ^ cout_1578; // @[Mul.scala 206:34]
  wire  cout_1678 = sum_1579 & cout_1578; // @[Mul.scala 207:34]
  wire  sum_1679 = sum_1580 ^ cout_1579; // @[Mul.scala 206:34]
  wire  sum_1698 = sum_1599 ^ cout_1598; // @[Mul.scala 206:34]
  wire  cout_1698 = sum_1599 & cout_1598; // @[Mul.scala 207:34]
  wire  sum_1699 = sum_1600 ^ cout_1599; // @[Mul.scala 206:34]
  wire  cout_1699 = sum_1600 & cout_1599; // @[Mul.scala 207:34]
  wire  sum_1700 = sum_1601 ^ cout_1600; // @[Mul.scala 206:34]
  wire  cout_1700 = sum_1601 & cout_1600; // @[Mul.scala 207:34]
  wire  _sum_T_2334 = sum_1602 ^ sum_1603; // @[Mul.scala 191:34]
  wire  sum_1701 = sum_1602 ^ sum_1603 ^ cout_1601; // @[Mul.scala 191:42]
  wire  cout_1701 = sum_1602 & sum_1603 | _sum_T_2334 & cout_1601; // @[Mul.scala 192:44]
  wire  sum_1702 = sum_1604 ^ sum_1605; // @[Mul.scala 206:34]
  wire  cout_1702 = sum_1604 & sum_1605; // @[Mul.scala 207:34]
  wire  sum_1703 = cout_1602 ^ cout_1603; // @[Mul.scala 206:34]
  wire  cout_1703 = cout_1602 & cout_1603; // @[Mul.scala 207:34]
  wire  sum_1704 = sum_1606 ^ sum_1607; // @[Mul.scala 206:34]
  wire  cout_1704 = sum_1606 & sum_1607; // @[Mul.scala 207:34]
  wire  sum_1705 = cout_1604 ^ cout_1605; // @[Mul.scala 206:34]
  wire  cout_1705 = cout_1604 & cout_1605; // @[Mul.scala 207:34]
  wire  sum_1706 = sum_1608 ^ sum_1609; // @[Mul.scala 206:34]
  wire  cout_1706 = sum_1608 & sum_1609; // @[Mul.scala 207:34]
  wire  sum_1707 = cout_1606 ^ cout_1607; // @[Mul.scala 206:34]
  wire  cout_1707 = cout_1606 & cout_1607; // @[Mul.scala 207:34]
  wire  sum_1708 = sum_1610 ^ sum_1611; // @[Mul.scala 206:34]
  wire  cout_1708 = sum_1610 & sum_1611; // @[Mul.scala 207:34]
  wire  sum_1709 = cout_1608 ^ cout_1609; // @[Mul.scala 206:34]
  wire  cout_1709 = cout_1608 & cout_1609; // @[Mul.scala 207:34]
  wire  sum_1710 = sum_1612 ^ sum_1613; // @[Mul.scala 206:34]
  wire  cout_1710 = sum_1612 & sum_1613; // @[Mul.scala 207:34]
  wire  sum_1711 = cout_1610 ^ cout_1611; // @[Mul.scala 206:34]
  wire  cout_1711 = cout_1610 & cout_1611; // @[Mul.scala 207:34]
  wire  sum_1712 = sum_1614 ^ sum_1615; // @[Mul.scala 206:34]
  wire  cout_1712 = sum_1614 & sum_1615; // @[Mul.scala 207:34]
  wire  sum_1713 = cout_1612 ^ cout_1613; // @[Mul.scala 206:34]
  wire  cout_1713 = cout_1612 & cout_1613; // @[Mul.scala 207:34]
  wire  sum_1714 = sum_1616 ^ sum_1617; // @[Mul.scala 206:34]
  wire  cout_1714 = sum_1616 & sum_1617; // @[Mul.scala 207:34]
  wire  sum_1715 = cout_1614 ^ cout_1615; // @[Mul.scala 206:34]
  wire  cout_1715 = cout_1614 & cout_1615; // @[Mul.scala 207:34]
  wire  sum_1716 = sum_1618 ^ sum_1619; // @[Mul.scala 206:34]
  wire  cout_1716 = sum_1618 & sum_1619; // @[Mul.scala 207:34]
  wire  sum_1717 = cout_1616 ^ cout_1617; // @[Mul.scala 206:34]
  wire  cout_1717 = cout_1616 & cout_1617; // @[Mul.scala 207:34]
  wire  sum_1718 = sum_1620 ^ sum_1621; // @[Mul.scala 206:34]
  wire  cout_1718 = sum_1620 & sum_1621; // @[Mul.scala 207:34]
  wire  sum_1719 = cout_1618 ^ cout_1619; // @[Mul.scala 206:34]
  wire  cout_1719 = cout_1618 & cout_1619; // @[Mul.scala 207:34]
  wire  sum_1720 = sum_1622 ^ sum_1623; // @[Mul.scala 206:34]
  wire  cout_1720 = sum_1622 & sum_1623; // @[Mul.scala 207:34]
  wire  sum_1721 = cout_1620 ^ cout_1621; // @[Mul.scala 206:34]
  wire  cout_1721 = cout_1620 & cout_1621; // @[Mul.scala 207:34]
  wire  sum_1722 = sum_1624 ^ sum_1625; // @[Mul.scala 206:34]
  wire  cout_1722 = sum_1624 & sum_1625; // @[Mul.scala 207:34]
  wire  sum_1723 = cout_1622 ^ cout_1623; // @[Mul.scala 206:34]
  wire  cout_1723 = cout_1622 & cout_1623; // @[Mul.scala 207:34]
  wire  sum_1724 = sum_1626 ^ sum_1627; // @[Mul.scala 206:34]
  wire  cout_1724 = sum_1626 & sum_1627; // @[Mul.scala 207:34]
  wire  sum_1725 = cout_1624 ^ cout_1625; // @[Mul.scala 206:34]
  wire  cout_1725 = cout_1624 & cout_1625; // @[Mul.scala 207:34]
  wire  sum_1726 = sum_1628 ^ sum_1629; // @[Mul.scala 206:34]
  wire  cout_1726 = sum_1628 & sum_1629; // @[Mul.scala 207:34]
  wire  sum_1727 = cout_1626 ^ cout_1627; // @[Mul.scala 206:34]
  wire  cout_1727 = cout_1626 & cout_1627; // @[Mul.scala 207:34]
  wire  sum_1728 = sum_1630 ^ sum_1631; // @[Mul.scala 206:34]
  wire  cout_1728 = sum_1630 & sum_1631; // @[Mul.scala 207:34]
  wire  sum_1729 = cout_1628 ^ cout_1629; // @[Mul.scala 206:34]
  wire  cout_1729 = cout_1628 & cout_1629; // @[Mul.scala 207:34]
  wire  sum_1730 = sum_1632 ^ sum_1633; // @[Mul.scala 206:34]
  wire  cout_1730 = sum_1632 & sum_1633; // @[Mul.scala 207:34]
  wire  sum_1731 = cout_1630 ^ cout_1631; // @[Mul.scala 206:34]
  wire  cout_1731 = cout_1630 & cout_1631; // @[Mul.scala 207:34]
  wire  sum_1732 = sum_1634 ^ sum_1635; // @[Mul.scala 206:34]
  wire  cout_1732 = sum_1634 & sum_1635; // @[Mul.scala 207:34]
  wire  sum_1733 = cout_1632 ^ cout_1633; // @[Mul.scala 206:34]
  wire  cout_1733 = cout_1632 & cout_1633; // @[Mul.scala 207:34]
  wire  sum_1734 = sum_1636 ^ sum_1637; // @[Mul.scala 206:34]
  wire  cout_1734 = sum_1636 & sum_1637; // @[Mul.scala 207:34]
  wire  sum_1735 = cout_1634 ^ cout_1635; // @[Mul.scala 206:34]
  wire  cout_1735 = cout_1634 & cout_1635; // @[Mul.scala 207:34]
  wire  sum_1736 = sum_1638 ^ sum_1639; // @[Mul.scala 206:34]
  wire  cout_1736 = sum_1638 & sum_1639; // @[Mul.scala 207:34]
  wire  sum_1737 = cout_1636 ^ cout_1637; // @[Mul.scala 206:34]
  wire  cout_1737 = cout_1636 & cout_1637; // @[Mul.scala 207:34]
  wire  sum_1738 = sum_1640 ^ sum_1641; // @[Mul.scala 206:34]
  wire  cout_1738 = sum_1640 & sum_1641; // @[Mul.scala 207:34]
  wire  sum_1739 = cout_1638 ^ cout_1639; // @[Mul.scala 206:34]
  wire  cout_1739 = cout_1638 & cout_1639; // @[Mul.scala 207:34]
  wire  sum_1740 = sum_1642 ^ sum_1643; // @[Mul.scala 206:34]
  wire  cout_1740 = sum_1642 & sum_1643; // @[Mul.scala 207:34]
  wire  sum_1741 = cout_1640 ^ cout_1641; // @[Mul.scala 206:34]
  wire  cout_1741 = cout_1640 & cout_1641; // @[Mul.scala 207:34]
  wire  sum_1742 = sum_1644 ^ sum_1645; // @[Mul.scala 206:34]
  wire  cout_1742 = sum_1644 & sum_1645; // @[Mul.scala 207:34]
  wire  sum_1743 = cout_1642 ^ cout_1643; // @[Mul.scala 206:34]
  wire  cout_1743 = cout_1642 & cout_1643; // @[Mul.scala 207:34]
  wire  sum_1744 = sum_1646 ^ sum_1647; // @[Mul.scala 206:34]
  wire  cout_1744 = sum_1646 & sum_1647; // @[Mul.scala 207:34]
  wire  sum_1745 = cout_1644 ^ cout_1645; // @[Mul.scala 206:34]
  wire  cout_1745 = cout_1644 & cout_1645; // @[Mul.scala 207:34]
  wire  sum_1746 = sum_1648 ^ sum_1649; // @[Mul.scala 206:34]
  wire  cout_1746 = sum_1648 & sum_1649; // @[Mul.scala 207:34]
  wire  sum_1747 = cout_1646 ^ cout_1647; // @[Mul.scala 206:34]
  wire  cout_1747 = cout_1646 & cout_1647; // @[Mul.scala 207:34]
  wire  sum_1748 = sum_1650 ^ sum_1651; // @[Mul.scala 206:34]
  wire  cout_1748 = sum_1650 & sum_1651; // @[Mul.scala 207:34]
  wire  sum_1749 = cout_1648 ^ cout_1649; // @[Mul.scala 206:34]
  wire  cout_1749 = cout_1648 & cout_1649; // @[Mul.scala 207:34]
  wire  sum_1750 = sum_1652 ^ sum_1653; // @[Mul.scala 206:34]
  wire  cout_1750 = sum_1652 & sum_1653; // @[Mul.scala 207:34]
  wire  sum_1751 = cout_1650 ^ cout_1651; // @[Mul.scala 206:34]
  wire  cout_1751 = cout_1650 & cout_1651; // @[Mul.scala 207:34]
  wire  sum_1752 = sum_1654 ^ sum_1655; // @[Mul.scala 206:34]
  wire  cout_1752 = sum_1654 & sum_1655; // @[Mul.scala 207:34]
  wire  sum_1753 = cout_1652 ^ cout_1653; // @[Mul.scala 206:34]
  wire  cout_1753 = cout_1652 & cout_1653; // @[Mul.scala 207:34]
  wire  sum_1754 = sum_1656 ^ sum_1657; // @[Mul.scala 206:34]
  wire  cout_1754 = sum_1656 & sum_1657; // @[Mul.scala 207:34]
  wire  sum_1755 = cout_1654 ^ cout_1655; // @[Mul.scala 206:34]
  wire  cout_1755 = cout_1654 & cout_1655; // @[Mul.scala 207:34]
  wire  sum_1756 = sum_1658 ^ sum_1659; // @[Mul.scala 206:34]
  wire  cout_1756 = sum_1658 & sum_1659; // @[Mul.scala 207:34]
  wire  sum_1757 = cout_1656 ^ cout_1657; // @[Mul.scala 206:34]
  wire  cout_1757 = cout_1656 & cout_1657; // @[Mul.scala 207:34]
  wire  sum_1758 = sum_1660 ^ sum_1661; // @[Mul.scala 206:34]
  wire  cout_1758 = sum_1660 & sum_1661; // @[Mul.scala 207:34]
  wire  sum_1759 = cout_1658 ^ cout_1659; // @[Mul.scala 206:34]
  wire  cout_1759 = cout_1658 & cout_1659; // @[Mul.scala 207:34]
  wire  sum_1760 = sum_1662 ^ sum_1663; // @[Mul.scala 206:34]
  wire  cout_1760 = sum_1662 & sum_1663; // @[Mul.scala 207:34]
  wire  sum_1761 = cout_1660 ^ cout_1661; // @[Mul.scala 206:34]
  wire  cout_1761 = cout_1660 & cout_1661; // @[Mul.scala 207:34]
  wire  sum_1762 = sum_1664 ^ sum_1665; // @[Mul.scala 206:34]
  wire  cout_1762 = sum_1664 & sum_1665; // @[Mul.scala 207:34]
  wire  sum_1763 = cout_1662 ^ cout_1663; // @[Mul.scala 206:34]
  wire  cout_1763 = cout_1662 & cout_1663; // @[Mul.scala 207:34]
  wire  sum_1764 = sum_1666 ^ sum_1667; // @[Mul.scala 206:34]
  wire  cout_1764 = sum_1666 & sum_1667; // @[Mul.scala 207:34]
  wire  sum_1765 = cout_1664 ^ cout_1665; // @[Mul.scala 206:34]
  wire  cout_1765 = cout_1664 & cout_1665; // @[Mul.scala 207:34]
  wire  sum_1766 = sum_1668 ^ sum_1669; // @[Mul.scala 206:34]
  wire  cout_1766 = sum_1668 & sum_1669; // @[Mul.scala 207:34]
  wire  sum_1767 = cout_1666 ^ cout_1667; // @[Mul.scala 206:34]
  wire  cout_1767 = cout_1666 & cout_1667; // @[Mul.scala 207:34]
  wire  sum_1768 = sum_1670 ^ sum_1671; // @[Mul.scala 206:34]
  wire  cout_1768 = sum_1670 & sum_1671; // @[Mul.scala 207:34]
  wire  sum_1769 = cout_1668 ^ cout_1669; // @[Mul.scala 206:34]
  wire  cout_1769 = cout_1668 & cout_1669; // @[Mul.scala 207:34]
  wire  sum_1770 = sum_1672 ^ sum_1673; // @[Mul.scala 206:34]
  wire  cout_1770 = sum_1672 & sum_1673; // @[Mul.scala 207:34]
  wire  sum_1771 = cout_1670 ^ cout_1671; // @[Mul.scala 206:34]
  wire  cout_1771 = cout_1670 & cout_1671; // @[Mul.scala 207:34]
  wire  _sum_T_2406 = sum_1674 ^ cout_1672; // @[Mul.scala 191:34]
  wire  sum_1772 = sum_1674 ^ cout_1672 ^ cout_1673; // @[Mul.scala 191:42]
  wire  cout_1772 = sum_1674 & cout_1672 | _sum_T_2406 & cout_1673; // @[Mul.scala 192:44]
  wire  sum_1773 = sum_1675 ^ cout_1674; // @[Mul.scala 206:34]
  wire  cout_1773 = sum_1675 & cout_1674; // @[Mul.scala 207:34]
  wire  sum_1774 = sum_1676 ^ cout_1675; // @[Mul.scala 206:34]
  wire  cout_1774 = sum_1676 & cout_1675; // @[Mul.scala 207:34]
  wire  sum_1775 = sum_1677 ^ cout_1676; // @[Mul.scala 206:34]
  wire  cout_1775 = sum_1677 & cout_1676; // @[Mul.scala 207:34]
  wire  sum_1776 = sum_1678 ^ cout_1677; // @[Mul.scala 206:34]
  wire  cout_1776 = sum_1678 & cout_1677; // @[Mul.scala 207:34]
  wire  sum_1777 = sum_1679 ^ cout_1678; // @[Mul.scala 206:34]
  wire  sum_1797 = sum_1699 ^ cout_1698; // @[Mul.scala 206:34]
  wire  cout_1797 = sum_1699 & cout_1698; // @[Mul.scala 207:34]
  wire  sum_1798 = sum_1700 ^ cout_1699; // @[Mul.scala 206:34]
  wire  cout_1798 = sum_1700 & cout_1699; // @[Mul.scala 207:34]
  wire  sum_1799 = sum_1701 ^ cout_1700; // @[Mul.scala 206:34]
  wire  cout_1799 = sum_1701 & cout_1700; // @[Mul.scala 207:34]
  wire  _sum_T_2435 = sum_1702 ^ sum_1703; // @[Mul.scala 191:34]
  wire  sum_1800 = sum_1702 ^ sum_1703 ^ cout_1701; // @[Mul.scala 191:42]
  wire  cout_1800 = sum_1702 & sum_1703 | _sum_T_2435 & cout_1701; // @[Mul.scala 192:44]
  wire  sum_1801 = sum_1704 ^ sum_1705; // @[Mul.scala 206:34]
  wire  cout_1801 = sum_1704 & sum_1705; // @[Mul.scala 207:34]
  wire  sum_1802 = cout_1702 ^ cout_1703; // @[Mul.scala 206:34]
  wire  cout_1802 = cout_1702 & cout_1703; // @[Mul.scala 207:34]
  wire  sum_1803 = sum_1706 ^ sum_1707; // @[Mul.scala 206:34]
  wire  cout_1803 = sum_1706 & sum_1707; // @[Mul.scala 207:34]
  wire  sum_1804 = cout_1704 ^ cout_1705; // @[Mul.scala 206:34]
  wire  cout_1804 = cout_1704 & cout_1705; // @[Mul.scala 207:34]
  wire  sum_1805 = sum_1708 ^ sum_1709; // @[Mul.scala 206:34]
  wire  cout_1805 = sum_1708 & sum_1709; // @[Mul.scala 207:34]
  wire  sum_1806 = cout_1706 ^ cout_1707; // @[Mul.scala 206:34]
  wire  cout_1806 = cout_1706 & cout_1707; // @[Mul.scala 207:34]
  wire  sum_1807 = sum_1710 ^ sum_1711; // @[Mul.scala 206:34]
  wire  cout_1807 = sum_1710 & sum_1711; // @[Mul.scala 207:34]
  wire  sum_1808 = cout_1708 ^ cout_1709; // @[Mul.scala 206:34]
  wire  cout_1808 = cout_1708 & cout_1709; // @[Mul.scala 207:34]
  wire  sum_1809 = sum_1712 ^ sum_1713; // @[Mul.scala 206:34]
  wire  cout_1809 = sum_1712 & sum_1713; // @[Mul.scala 207:34]
  wire  sum_1810 = cout_1710 ^ cout_1711; // @[Mul.scala 206:34]
  wire  cout_1810 = cout_1710 & cout_1711; // @[Mul.scala 207:34]
  wire  sum_1811 = sum_1714 ^ sum_1715; // @[Mul.scala 206:34]
  wire  cout_1811 = sum_1714 & sum_1715; // @[Mul.scala 207:34]
  wire  sum_1812 = cout_1712 ^ cout_1713; // @[Mul.scala 206:34]
  wire  cout_1812 = cout_1712 & cout_1713; // @[Mul.scala 207:34]
  wire  sum_1813 = sum_1716 ^ sum_1717; // @[Mul.scala 206:34]
  wire  cout_1813 = sum_1716 & sum_1717; // @[Mul.scala 207:34]
  wire  sum_1814 = cout_1714 ^ cout_1715; // @[Mul.scala 206:34]
  wire  cout_1814 = cout_1714 & cout_1715; // @[Mul.scala 207:34]
  wire  sum_1815 = sum_1718 ^ sum_1719; // @[Mul.scala 206:34]
  wire  cout_1815 = sum_1718 & sum_1719; // @[Mul.scala 207:34]
  wire  sum_1816 = cout_1716 ^ cout_1717; // @[Mul.scala 206:34]
  wire  cout_1816 = cout_1716 & cout_1717; // @[Mul.scala 207:34]
  wire  sum_1817 = sum_1720 ^ sum_1721; // @[Mul.scala 206:34]
  wire  cout_1817 = sum_1720 & sum_1721; // @[Mul.scala 207:34]
  wire  sum_1818 = cout_1718 ^ cout_1719; // @[Mul.scala 206:34]
  wire  cout_1818 = cout_1718 & cout_1719; // @[Mul.scala 207:34]
  wire  sum_1819 = sum_1722 ^ sum_1723; // @[Mul.scala 206:34]
  wire  cout_1819 = sum_1722 & sum_1723; // @[Mul.scala 207:34]
  wire  sum_1820 = cout_1720 ^ cout_1721; // @[Mul.scala 206:34]
  wire  cout_1820 = cout_1720 & cout_1721; // @[Mul.scala 207:34]
  wire  sum_1821 = sum_1724 ^ sum_1725; // @[Mul.scala 206:34]
  wire  cout_1821 = sum_1724 & sum_1725; // @[Mul.scala 207:34]
  wire  sum_1822 = cout_1722 ^ cout_1723; // @[Mul.scala 206:34]
  wire  cout_1822 = cout_1722 & cout_1723; // @[Mul.scala 207:34]
  wire  sum_1823 = sum_1726 ^ sum_1727; // @[Mul.scala 206:34]
  wire  cout_1823 = sum_1726 & sum_1727; // @[Mul.scala 207:34]
  wire  sum_1824 = cout_1724 ^ cout_1725; // @[Mul.scala 206:34]
  wire  cout_1824 = cout_1724 & cout_1725; // @[Mul.scala 207:34]
  wire  sum_1825 = sum_1728 ^ sum_1729; // @[Mul.scala 206:34]
  wire  cout_1825 = sum_1728 & sum_1729; // @[Mul.scala 207:34]
  wire  sum_1826 = cout_1726 ^ cout_1727; // @[Mul.scala 206:34]
  wire  cout_1826 = cout_1726 & cout_1727; // @[Mul.scala 207:34]
  wire  sum_1827 = sum_1730 ^ sum_1731; // @[Mul.scala 206:34]
  wire  cout_1827 = sum_1730 & sum_1731; // @[Mul.scala 207:34]
  wire  sum_1828 = cout_1728 ^ cout_1729; // @[Mul.scala 206:34]
  wire  cout_1828 = cout_1728 & cout_1729; // @[Mul.scala 207:34]
  wire  sum_1829 = sum_1732 ^ sum_1733; // @[Mul.scala 206:34]
  wire  cout_1829 = sum_1732 & sum_1733; // @[Mul.scala 207:34]
  wire  sum_1830 = cout_1730 ^ cout_1731; // @[Mul.scala 206:34]
  wire  cout_1830 = cout_1730 & cout_1731; // @[Mul.scala 207:34]
  wire  sum_1831 = sum_1734 ^ sum_1735; // @[Mul.scala 206:34]
  wire  cout_1831 = sum_1734 & sum_1735; // @[Mul.scala 207:34]
  wire  sum_1832 = cout_1732 ^ cout_1733; // @[Mul.scala 206:34]
  wire  cout_1832 = cout_1732 & cout_1733; // @[Mul.scala 207:34]
  wire  sum_1833 = sum_1736 ^ sum_1737; // @[Mul.scala 206:34]
  wire  cout_1833 = sum_1736 & sum_1737; // @[Mul.scala 207:34]
  wire  sum_1834 = cout_1734 ^ cout_1735; // @[Mul.scala 206:34]
  wire  cout_1834 = cout_1734 & cout_1735; // @[Mul.scala 207:34]
  wire  sum_1835 = sum_1738 ^ sum_1739; // @[Mul.scala 206:34]
  wire  cout_1835 = sum_1738 & sum_1739; // @[Mul.scala 207:34]
  wire  sum_1836 = cout_1736 ^ cout_1737; // @[Mul.scala 206:34]
  wire  cout_1836 = cout_1736 & cout_1737; // @[Mul.scala 207:34]
  wire  sum_1837 = sum_1740 ^ sum_1741; // @[Mul.scala 206:34]
  wire  cout_1837 = sum_1740 & sum_1741; // @[Mul.scala 207:34]
  wire  sum_1838 = cout_1738 ^ cout_1739; // @[Mul.scala 206:34]
  wire  cout_1838 = cout_1738 & cout_1739; // @[Mul.scala 207:34]
  wire  sum_1839 = sum_1742 ^ sum_1743; // @[Mul.scala 206:34]
  wire  cout_1839 = sum_1742 & sum_1743; // @[Mul.scala 207:34]
  wire  sum_1840 = cout_1740 ^ cout_1741; // @[Mul.scala 206:34]
  wire  cout_1840 = cout_1740 & cout_1741; // @[Mul.scala 207:34]
  wire  sum_1841 = sum_1744 ^ sum_1745; // @[Mul.scala 206:34]
  wire  cout_1841 = sum_1744 & sum_1745; // @[Mul.scala 207:34]
  wire  sum_1842 = cout_1742 ^ cout_1743; // @[Mul.scala 206:34]
  wire  cout_1842 = cout_1742 & cout_1743; // @[Mul.scala 207:34]
  wire  sum_1843 = sum_1746 ^ sum_1747; // @[Mul.scala 206:34]
  wire  cout_1843 = sum_1746 & sum_1747; // @[Mul.scala 207:34]
  wire  sum_1844 = cout_1744 ^ cout_1745; // @[Mul.scala 206:34]
  wire  cout_1844 = cout_1744 & cout_1745; // @[Mul.scala 207:34]
  wire  sum_1845 = sum_1748 ^ sum_1749; // @[Mul.scala 206:34]
  wire  cout_1845 = sum_1748 & sum_1749; // @[Mul.scala 207:34]
  wire  sum_1846 = cout_1746 ^ cout_1747; // @[Mul.scala 206:34]
  wire  cout_1846 = cout_1746 & cout_1747; // @[Mul.scala 207:34]
  wire  sum_1847 = sum_1750 ^ sum_1751; // @[Mul.scala 206:34]
  wire  cout_1847 = sum_1750 & sum_1751; // @[Mul.scala 207:34]
  wire  sum_1848 = cout_1748 ^ cout_1749; // @[Mul.scala 206:34]
  wire  cout_1848 = cout_1748 & cout_1749; // @[Mul.scala 207:34]
  wire  sum_1849 = sum_1752 ^ sum_1753; // @[Mul.scala 206:34]
  wire  cout_1849 = sum_1752 & sum_1753; // @[Mul.scala 207:34]
  wire  sum_1850 = cout_1750 ^ cout_1751; // @[Mul.scala 206:34]
  wire  cout_1850 = cout_1750 & cout_1751; // @[Mul.scala 207:34]
  wire  sum_1851 = sum_1754 ^ sum_1755; // @[Mul.scala 206:34]
  wire  cout_1851 = sum_1754 & sum_1755; // @[Mul.scala 207:34]
  wire  sum_1852 = cout_1752 ^ cout_1753; // @[Mul.scala 206:34]
  wire  cout_1852 = cout_1752 & cout_1753; // @[Mul.scala 207:34]
  wire  sum_1853 = sum_1756 ^ sum_1757; // @[Mul.scala 206:34]
  wire  cout_1853 = sum_1756 & sum_1757; // @[Mul.scala 207:34]
  wire  sum_1854 = cout_1754 ^ cout_1755; // @[Mul.scala 206:34]
  wire  cout_1854 = cout_1754 & cout_1755; // @[Mul.scala 207:34]
  wire  sum_1855 = sum_1758 ^ sum_1759; // @[Mul.scala 206:34]
  wire  cout_1855 = sum_1758 & sum_1759; // @[Mul.scala 207:34]
  wire  sum_1856 = cout_1756 ^ cout_1757; // @[Mul.scala 206:34]
  wire  cout_1856 = cout_1756 & cout_1757; // @[Mul.scala 207:34]
  wire  sum_1857 = sum_1760 ^ sum_1761; // @[Mul.scala 206:34]
  wire  cout_1857 = sum_1760 & sum_1761; // @[Mul.scala 207:34]
  wire  sum_1858 = cout_1758 ^ cout_1759; // @[Mul.scala 206:34]
  wire  cout_1858 = cout_1758 & cout_1759; // @[Mul.scala 207:34]
  wire  sum_1859 = sum_1762 ^ sum_1763; // @[Mul.scala 206:34]
  wire  cout_1859 = sum_1762 & sum_1763; // @[Mul.scala 207:34]
  wire  sum_1860 = cout_1760 ^ cout_1761; // @[Mul.scala 206:34]
  wire  cout_1860 = cout_1760 & cout_1761; // @[Mul.scala 207:34]
  wire  sum_1861 = sum_1764 ^ sum_1765; // @[Mul.scala 206:34]
  wire  cout_1861 = sum_1764 & sum_1765; // @[Mul.scala 207:34]
  wire  sum_1862 = cout_1762 ^ cout_1763; // @[Mul.scala 206:34]
  wire  cout_1862 = cout_1762 & cout_1763; // @[Mul.scala 207:34]
  wire  sum_1863 = sum_1766 ^ sum_1767; // @[Mul.scala 206:34]
  wire  cout_1863 = sum_1766 & sum_1767; // @[Mul.scala 207:34]
  wire  sum_1864 = cout_1764 ^ cout_1765; // @[Mul.scala 206:34]
  wire  cout_1864 = cout_1764 & cout_1765; // @[Mul.scala 207:34]
  wire  sum_1865 = sum_1768 ^ sum_1769; // @[Mul.scala 206:34]
  wire  cout_1865 = sum_1768 & sum_1769; // @[Mul.scala 207:34]
  wire  sum_1866 = cout_1766 ^ cout_1767; // @[Mul.scala 206:34]
  wire  cout_1866 = cout_1766 & cout_1767; // @[Mul.scala 207:34]
  wire  sum_1867 = sum_1770 ^ sum_1771; // @[Mul.scala 206:34]
  wire  cout_1867 = sum_1770 & sum_1771; // @[Mul.scala 207:34]
  wire  sum_1868 = cout_1768 ^ cout_1769; // @[Mul.scala 206:34]
  wire  cout_1868 = cout_1768 & cout_1769; // @[Mul.scala 207:34]
  wire  _sum_T_2505 = sum_1772 ^ cout_1770; // @[Mul.scala 191:34]
  wire  sum_1869 = sum_1772 ^ cout_1770 ^ cout_1771; // @[Mul.scala 191:42]
  wire  cout_1869 = sum_1772 & cout_1770 | _sum_T_2505 & cout_1771; // @[Mul.scala 192:44]
  wire  sum_1870 = sum_1773 ^ cout_1772; // @[Mul.scala 206:34]
  wire  cout_1870 = sum_1773 & cout_1772; // @[Mul.scala 207:34]
  wire  sum_1871 = sum_1774 ^ cout_1773; // @[Mul.scala 206:34]
  wire  cout_1871 = sum_1774 & cout_1773; // @[Mul.scala 207:34]
  wire  sum_1872 = sum_1775 ^ cout_1774; // @[Mul.scala 206:34]
  wire  cout_1872 = sum_1775 & cout_1774; // @[Mul.scala 207:34]
  wire  sum_1873 = sum_1776 ^ cout_1775; // @[Mul.scala 206:34]
  wire  cout_1873 = sum_1776 & cout_1775; // @[Mul.scala 207:34]
  wire  sum_1874 = sum_1777 ^ cout_1776; // @[Mul.scala 206:34]
  wire  sum_1895 = sum_1798 ^ cout_1797; // @[Mul.scala 206:34]
  wire  cout_1895 = sum_1798 & cout_1797; // @[Mul.scala 207:34]
  wire  sum_1896 = sum_1799 ^ cout_1798; // @[Mul.scala 206:34]
  wire  cout_1896 = sum_1799 & cout_1798; // @[Mul.scala 207:34]
  wire  sum_1897 = sum_1800 ^ cout_1799; // @[Mul.scala 206:34]
  wire  cout_1897 = sum_1800 & cout_1799; // @[Mul.scala 207:34]
  wire  _sum_T_2535 = sum_1801 ^ sum_1802; // @[Mul.scala 191:34]
  wire  sum_1898 = sum_1801 ^ sum_1802 ^ cout_1800; // @[Mul.scala 191:42]
  wire  cout_1898 = sum_1801 & sum_1802 | _sum_T_2535 & cout_1800; // @[Mul.scala 192:44]
  wire  sum_1899 = sum_1803 ^ sum_1804; // @[Mul.scala 206:34]
  wire  cout_1899 = sum_1803 & sum_1804; // @[Mul.scala 207:34]
  wire  sum_1900 = cout_1801 ^ cout_1802; // @[Mul.scala 206:34]
  wire  cout_1900 = cout_1801 & cout_1802; // @[Mul.scala 207:34]
  wire  sum_1901 = sum_1805 ^ sum_1806; // @[Mul.scala 206:34]
  wire  cout_1901 = sum_1805 & sum_1806; // @[Mul.scala 207:34]
  wire  sum_1902 = cout_1803 ^ cout_1804; // @[Mul.scala 206:34]
  wire  cout_1902 = cout_1803 & cout_1804; // @[Mul.scala 207:34]
  wire  sum_1903 = sum_1807 ^ sum_1808; // @[Mul.scala 206:34]
  wire  cout_1903 = sum_1807 & sum_1808; // @[Mul.scala 207:34]
  wire  sum_1904 = cout_1805 ^ cout_1806; // @[Mul.scala 206:34]
  wire  cout_1904 = cout_1805 & cout_1806; // @[Mul.scala 207:34]
  wire  sum_1905 = sum_1809 ^ sum_1810; // @[Mul.scala 206:34]
  wire  cout_1905 = sum_1809 & sum_1810; // @[Mul.scala 207:34]
  wire  sum_1906 = cout_1807 ^ cout_1808; // @[Mul.scala 206:34]
  wire  cout_1906 = cout_1807 & cout_1808; // @[Mul.scala 207:34]
  wire  sum_1907 = sum_1811 ^ sum_1812; // @[Mul.scala 206:34]
  wire  cout_1907 = sum_1811 & sum_1812; // @[Mul.scala 207:34]
  wire  sum_1908 = cout_1809 ^ cout_1810; // @[Mul.scala 206:34]
  wire  cout_1908 = cout_1809 & cout_1810; // @[Mul.scala 207:34]
  wire  sum_1909 = sum_1813 ^ sum_1814; // @[Mul.scala 206:34]
  wire  cout_1909 = sum_1813 & sum_1814; // @[Mul.scala 207:34]
  wire  sum_1910 = cout_1811 ^ cout_1812; // @[Mul.scala 206:34]
  wire  cout_1910 = cout_1811 & cout_1812; // @[Mul.scala 207:34]
  wire  sum_1911 = sum_1815 ^ sum_1816; // @[Mul.scala 206:34]
  wire  cout_1911 = sum_1815 & sum_1816; // @[Mul.scala 207:34]
  wire  sum_1912 = cout_1813 ^ cout_1814; // @[Mul.scala 206:34]
  wire  cout_1912 = cout_1813 & cout_1814; // @[Mul.scala 207:34]
  wire  sum_1913 = sum_1817 ^ sum_1818; // @[Mul.scala 206:34]
  wire  cout_1913 = sum_1817 & sum_1818; // @[Mul.scala 207:34]
  wire  sum_1914 = cout_1815 ^ cout_1816; // @[Mul.scala 206:34]
  wire  cout_1914 = cout_1815 & cout_1816; // @[Mul.scala 207:34]
  wire  sum_1915 = sum_1819 ^ sum_1820; // @[Mul.scala 206:34]
  wire  cout_1915 = sum_1819 & sum_1820; // @[Mul.scala 207:34]
  wire  sum_1916 = cout_1817 ^ cout_1818; // @[Mul.scala 206:34]
  wire  cout_1916 = cout_1817 & cout_1818; // @[Mul.scala 207:34]
  wire  sum_1917 = sum_1821 ^ sum_1822; // @[Mul.scala 206:34]
  wire  cout_1917 = sum_1821 & sum_1822; // @[Mul.scala 207:34]
  wire  sum_1918 = cout_1819 ^ cout_1820; // @[Mul.scala 206:34]
  wire  cout_1918 = cout_1819 & cout_1820; // @[Mul.scala 207:34]
  wire  sum_1919 = sum_1823 ^ sum_1824; // @[Mul.scala 206:34]
  wire  cout_1919 = sum_1823 & sum_1824; // @[Mul.scala 207:34]
  wire  sum_1920 = cout_1821 ^ cout_1822; // @[Mul.scala 206:34]
  wire  cout_1920 = cout_1821 & cout_1822; // @[Mul.scala 207:34]
  wire  sum_1921 = sum_1825 ^ sum_1826; // @[Mul.scala 206:34]
  wire  cout_1921 = sum_1825 & sum_1826; // @[Mul.scala 207:34]
  wire  sum_1922 = cout_1823 ^ cout_1824; // @[Mul.scala 206:34]
  wire  cout_1922 = cout_1823 & cout_1824; // @[Mul.scala 207:34]
  wire  sum_1923 = sum_1827 ^ sum_1828; // @[Mul.scala 206:34]
  wire  cout_1923 = sum_1827 & sum_1828; // @[Mul.scala 207:34]
  wire  sum_1924 = cout_1825 ^ cout_1826; // @[Mul.scala 206:34]
  wire  cout_1924 = cout_1825 & cout_1826; // @[Mul.scala 207:34]
  wire  sum_1925 = sum_1829 ^ sum_1830; // @[Mul.scala 206:34]
  wire  cout_1925 = sum_1829 & sum_1830; // @[Mul.scala 207:34]
  wire  sum_1926 = cout_1827 ^ cout_1828; // @[Mul.scala 206:34]
  wire  cout_1926 = cout_1827 & cout_1828; // @[Mul.scala 207:34]
  wire  sum_1927 = sum_1831 ^ sum_1832; // @[Mul.scala 206:34]
  wire  cout_1927 = sum_1831 & sum_1832; // @[Mul.scala 207:34]
  wire  sum_1928 = cout_1829 ^ cout_1830; // @[Mul.scala 206:34]
  wire  cout_1928 = cout_1829 & cout_1830; // @[Mul.scala 207:34]
  wire  sum_1929 = sum_1833 ^ sum_1834; // @[Mul.scala 206:34]
  wire  cout_1929 = sum_1833 & sum_1834; // @[Mul.scala 207:34]
  wire  sum_1930 = cout_1831 ^ cout_1832; // @[Mul.scala 206:34]
  wire  cout_1930 = cout_1831 & cout_1832; // @[Mul.scala 207:34]
  wire  sum_1931 = sum_1835 ^ sum_1836; // @[Mul.scala 206:34]
  wire  cout_1931 = sum_1835 & sum_1836; // @[Mul.scala 207:34]
  wire  sum_1932 = cout_1833 ^ cout_1834; // @[Mul.scala 206:34]
  wire  cout_1932 = cout_1833 & cout_1834; // @[Mul.scala 207:34]
  wire  sum_1933 = sum_1837 ^ sum_1838; // @[Mul.scala 206:34]
  wire  cout_1933 = sum_1837 & sum_1838; // @[Mul.scala 207:34]
  wire  sum_1934 = cout_1835 ^ cout_1836; // @[Mul.scala 206:34]
  wire  cout_1934 = cout_1835 & cout_1836; // @[Mul.scala 207:34]
  wire  sum_1935 = sum_1839 ^ sum_1840; // @[Mul.scala 206:34]
  wire  cout_1935 = sum_1839 & sum_1840; // @[Mul.scala 207:34]
  wire  sum_1936 = cout_1837 ^ cout_1838; // @[Mul.scala 206:34]
  wire  cout_1936 = cout_1837 & cout_1838; // @[Mul.scala 207:34]
  wire  sum_1937 = sum_1841 ^ sum_1842; // @[Mul.scala 206:34]
  wire  cout_1937 = sum_1841 & sum_1842; // @[Mul.scala 207:34]
  wire  sum_1938 = cout_1839 ^ cout_1840; // @[Mul.scala 206:34]
  wire  cout_1938 = cout_1839 & cout_1840; // @[Mul.scala 207:34]
  wire  sum_1939 = sum_1843 ^ sum_1844; // @[Mul.scala 206:34]
  wire  cout_1939 = sum_1843 & sum_1844; // @[Mul.scala 207:34]
  wire  sum_1940 = cout_1841 ^ cout_1842; // @[Mul.scala 206:34]
  wire  cout_1940 = cout_1841 & cout_1842; // @[Mul.scala 207:34]
  wire  sum_1941 = sum_1845 ^ sum_1846; // @[Mul.scala 206:34]
  wire  cout_1941 = sum_1845 & sum_1846; // @[Mul.scala 207:34]
  wire  sum_1942 = cout_1843 ^ cout_1844; // @[Mul.scala 206:34]
  wire  cout_1942 = cout_1843 & cout_1844; // @[Mul.scala 207:34]
  wire  sum_1943 = sum_1847 ^ sum_1848; // @[Mul.scala 206:34]
  wire  cout_1943 = sum_1847 & sum_1848; // @[Mul.scala 207:34]
  wire  sum_1944 = cout_1845 ^ cout_1846; // @[Mul.scala 206:34]
  wire  cout_1944 = cout_1845 & cout_1846; // @[Mul.scala 207:34]
  wire  sum_1945 = sum_1849 ^ sum_1850; // @[Mul.scala 206:34]
  wire  cout_1945 = sum_1849 & sum_1850; // @[Mul.scala 207:34]
  wire  sum_1946 = cout_1847 ^ cout_1848; // @[Mul.scala 206:34]
  wire  cout_1946 = cout_1847 & cout_1848; // @[Mul.scala 207:34]
  wire  sum_1947 = sum_1851 ^ sum_1852; // @[Mul.scala 206:34]
  wire  cout_1947 = sum_1851 & sum_1852; // @[Mul.scala 207:34]
  wire  sum_1948 = cout_1849 ^ cout_1850; // @[Mul.scala 206:34]
  wire  cout_1948 = cout_1849 & cout_1850; // @[Mul.scala 207:34]
  wire  sum_1949 = sum_1853 ^ sum_1854; // @[Mul.scala 206:34]
  wire  cout_1949 = sum_1853 & sum_1854; // @[Mul.scala 207:34]
  wire  sum_1950 = cout_1851 ^ cout_1852; // @[Mul.scala 206:34]
  wire  cout_1950 = cout_1851 & cout_1852; // @[Mul.scala 207:34]
  wire  sum_1951 = sum_1855 ^ sum_1856; // @[Mul.scala 206:34]
  wire  cout_1951 = sum_1855 & sum_1856; // @[Mul.scala 207:34]
  wire  sum_1952 = cout_1853 ^ cout_1854; // @[Mul.scala 206:34]
  wire  cout_1952 = cout_1853 & cout_1854; // @[Mul.scala 207:34]
  wire  sum_1953 = sum_1857 ^ sum_1858; // @[Mul.scala 206:34]
  wire  cout_1953 = sum_1857 & sum_1858; // @[Mul.scala 207:34]
  wire  sum_1954 = cout_1855 ^ cout_1856; // @[Mul.scala 206:34]
  wire  cout_1954 = cout_1855 & cout_1856; // @[Mul.scala 207:34]
  wire  sum_1955 = sum_1859 ^ sum_1860; // @[Mul.scala 206:34]
  wire  cout_1955 = sum_1859 & sum_1860; // @[Mul.scala 207:34]
  wire  sum_1956 = cout_1857 ^ cout_1858; // @[Mul.scala 206:34]
  wire  cout_1956 = cout_1857 & cout_1858; // @[Mul.scala 207:34]
  wire  sum_1957 = sum_1861 ^ sum_1862; // @[Mul.scala 206:34]
  wire  cout_1957 = sum_1861 & sum_1862; // @[Mul.scala 207:34]
  wire  sum_1958 = cout_1859 ^ cout_1860; // @[Mul.scala 206:34]
  wire  cout_1958 = cout_1859 & cout_1860; // @[Mul.scala 207:34]
  wire  sum_1959 = sum_1863 ^ sum_1864; // @[Mul.scala 206:34]
  wire  cout_1959 = sum_1863 & sum_1864; // @[Mul.scala 207:34]
  wire  sum_1960 = cout_1861 ^ cout_1862; // @[Mul.scala 206:34]
  wire  cout_1960 = cout_1861 & cout_1862; // @[Mul.scala 207:34]
  wire  sum_1961 = sum_1865 ^ sum_1866; // @[Mul.scala 206:34]
  wire  cout_1961 = sum_1865 & sum_1866; // @[Mul.scala 207:34]
  wire  sum_1962 = cout_1863 ^ cout_1864; // @[Mul.scala 206:34]
  wire  cout_1962 = cout_1863 & cout_1864; // @[Mul.scala 207:34]
  wire  sum_1963 = sum_1867 ^ sum_1868; // @[Mul.scala 206:34]
  wire  cout_1963 = sum_1867 & sum_1868; // @[Mul.scala 207:34]
  wire  sum_1964 = cout_1865 ^ cout_1866; // @[Mul.scala 206:34]
  wire  cout_1964 = cout_1865 & cout_1866; // @[Mul.scala 207:34]
  wire  _sum_T_2603 = sum_1869 ^ cout_1867; // @[Mul.scala 191:34]
  wire  sum_1965 = sum_1869 ^ cout_1867 ^ cout_1868; // @[Mul.scala 191:42]
  wire  cout_1965 = sum_1869 & cout_1867 | _sum_T_2603 & cout_1868; // @[Mul.scala 192:44]
  wire  sum_1966 = sum_1870 ^ cout_1869; // @[Mul.scala 206:34]
  wire  cout_1966 = sum_1870 & cout_1869; // @[Mul.scala 207:34]
  wire  sum_1967 = sum_1871 ^ cout_1870; // @[Mul.scala 206:34]
  wire  cout_1967 = sum_1871 & cout_1870; // @[Mul.scala 207:34]
  wire  sum_1968 = sum_1872 ^ cout_1871; // @[Mul.scala 206:34]
  wire  cout_1968 = sum_1872 & cout_1871; // @[Mul.scala 207:34]
  wire  sum_1969 = sum_1873 ^ cout_1872; // @[Mul.scala 206:34]
  wire  cout_1969 = sum_1873 & cout_1872; // @[Mul.scala 207:34]
  wire  sum_1970 = sum_1874 ^ cout_1873; // @[Mul.scala 206:34]
  wire  sum_1992 = sum_1896 ^ cout_1895; // @[Mul.scala 206:34]
  wire  cout_1992 = sum_1896 & cout_1895; // @[Mul.scala 207:34]
  wire  sum_1993 = sum_1897 ^ cout_1896; // @[Mul.scala 206:34]
  wire  cout_1993 = sum_1897 & cout_1896; // @[Mul.scala 207:34]
  wire  sum_1994 = sum_1898 ^ cout_1897; // @[Mul.scala 206:34]
  wire  cout_1994 = sum_1898 & cout_1897; // @[Mul.scala 207:34]
  wire  _sum_T_2634 = sum_1899 ^ sum_1900; // @[Mul.scala 191:34]
  wire  sum_1995 = sum_1899 ^ sum_1900 ^ cout_1898; // @[Mul.scala 191:42]
  wire  cout_1995 = sum_1899 & sum_1900 | _sum_T_2634 & cout_1898; // @[Mul.scala 192:44]
  wire  sum_1996 = sum_1901 ^ sum_1902; // @[Mul.scala 206:34]
  wire  cout_1996 = sum_1901 & sum_1902; // @[Mul.scala 207:34]
  wire  sum_1997 = cout_1899 ^ cout_1900; // @[Mul.scala 206:34]
  wire  cout_1997 = cout_1899 & cout_1900; // @[Mul.scala 207:34]
  wire  sum_1998 = sum_1903 ^ sum_1904; // @[Mul.scala 206:34]
  wire  cout_1998 = sum_1903 & sum_1904; // @[Mul.scala 207:34]
  wire  sum_1999 = cout_1901 ^ cout_1902; // @[Mul.scala 206:34]
  wire  cout_1999 = cout_1901 & cout_1902; // @[Mul.scala 207:34]
  wire  sum_2000 = sum_1905 ^ sum_1906; // @[Mul.scala 206:34]
  wire  cout_2000 = sum_1905 & sum_1906; // @[Mul.scala 207:34]
  wire  sum_2001 = cout_1903 ^ cout_1904; // @[Mul.scala 206:34]
  wire  cout_2001 = cout_1903 & cout_1904; // @[Mul.scala 207:34]
  wire  sum_2002 = sum_1907 ^ sum_1908; // @[Mul.scala 206:34]
  wire  cout_2002 = sum_1907 & sum_1908; // @[Mul.scala 207:34]
  wire  sum_2003 = cout_1905 ^ cout_1906; // @[Mul.scala 206:34]
  wire  cout_2003 = cout_1905 & cout_1906; // @[Mul.scala 207:34]
  wire  sum_2004 = sum_1909 ^ sum_1910; // @[Mul.scala 206:34]
  wire  cout_2004 = sum_1909 & sum_1910; // @[Mul.scala 207:34]
  wire  sum_2005 = cout_1907 ^ cout_1908; // @[Mul.scala 206:34]
  wire  cout_2005 = cout_1907 & cout_1908; // @[Mul.scala 207:34]
  wire  sum_2006 = sum_1911 ^ sum_1912; // @[Mul.scala 206:34]
  wire  cout_2006 = sum_1911 & sum_1912; // @[Mul.scala 207:34]
  wire  sum_2007 = cout_1909 ^ cout_1910; // @[Mul.scala 206:34]
  wire  cout_2007 = cout_1909 & cout_1910; // @[Mul.scala 207:34]
  wire  sum_2008 = sum_1913 ^ sum_1914; // @[Mul.scala 206:34]
  wire  cout_2008 = sum_1913 & sum_1914; // @[Mul.scala 207:34]
  wire  sum_2009 = cout_1911 ^ cout_1912; // @[Mul.scala 206:34]
  wire  cout_2009 = cout_1911 & cout_1912; // @[Mul.scala 207:34]
  wire  sum_2010 = sum_1915 ^ sum_1916; // @[Mul.scala 206:34]
  wire  cout_2010 = sum_1915 & sum_1916; // @[Mul.scala 207:34]
  wire  sum_2011 = cout_1913 ^ cout_1914; // @[Mul.scala 206:34]
  wire  cout_2011 = cout_1913 & cout_1914; // @[Mul.scala 207:34]
  wire  sum_2012 = sum_1917 ^ sum_1918; // @[Mul.scala 206:34]
  wire  cout_2012 = sum_1917 & sum_1918; // @[Mul.scala 207:34]
  wire  sum_2013 = cout_1915 ^ cout_1916; // @[Mul.scala 206:34]
  wire  cout_2013 = cout_1915 & cout_1916; // @[Mul.scala 207:34]
  wire  sum_2014 = sum_1919 ^ sum_1920; // @[Mul.scala 206:34]
  wire  cout_2014 = sum_1919 & sum_1920; // @[Mul.scala 207:34]
  wire  sum_2015 = cout_1917 ^ cout_1918; // @[Mul.scala 206:34]
  wire  cout_2015 = cout_1917 & cout_1918; // @[Mul.scala 207:34]
  wire  sum_2016 = sum_1921 ^ sum_1922; // @[Mul.scala 206:34]
  wire  cout_2016 = sum_1921 & sum_1922; // @[Mul.scala 207:34]
  wire  sum_2017 = cout_1919 ^ cout_1920; // @[Mul.scala 206:34]
  wire  cout_2017 = cout_1919 & cout_1920; // @[Mul.scala 207:34]
  wire  sum_2018 = sum_1923 ^ sum_1924; // @[Mul.scala 206:34]
  wire  cout_2018 = sum_1923 & sum_1924; // @[Mul.scala 207:34]
  wire  sum_2019 = cout_1921 ^ cout_1922; // @[Mul.scala 206:34]
  wire  cout_2019 = cout_1921 & cout_1922; // @[Mul.scala 207:34]
  wire  sum_2020 = sum_1925 ^ sum_1926; // @[Mul.scala 206:34]
  wire  cout_2020 = sum_1925 & sum_1926; // @[Mul.scala 207:34]
  wire  sum_2021 = cout_1923 ^ cout_1924; // @[Mul.scala 206:34]
  wire  cout_2021 = cout_1923 & cout_1924; // @[Mul.scala 207:34]
  wire  sum_2022 = sum_1927 ^ sum_1928; // @[Mul.scala 206:34]
  wire  cout_2022 = sum_1927 & sum_1928; // @[Mul.scala 207:34]
  wire  sum_2023 = cout_1925 ^ cout_1926; // @[Mul.scala 206:34]
  wire  cout_2023 = cout_1925 & cout_1926; // @[Mul.scala 207:34]
  wire  sum_2024 = sum_1929 ^ sum_1930; // @[Mul.scala 206:34]
  wire  cout_2024 = sum_1929 & sum_1930; // @[Mul.scala 207:34]
  wire  sum_2025 = cout_1927 ^ cout_1928; // @[Mul.scala 206:34]
  wire  cout_2025 = cout_1927 & cout_1928; // @[Mul.scala 207:34]
  wire  sum_2026 = sum_1931 ^ sum_1932; // @[Mul.scala 206:34]
  wire  cout_2026 = sum_1931 & sum_1932; // @[Mul.scala 207:34]
  wire  sum_2027 = cout_1929 ^ cout_1930; // @[Mul.scala 206:34]
  wire  cout_2027 = cout_1929 & cout_1930; // @[Mul.scala 207:34]
  wire  sum_2028 = sum_1933 ^ sum_1934; // @[Mul.scala 206:34]
  wire  cout_2028 = sum_1933 & sum_1934; // @[Mul.scala 207:34]
  wire  sum_2029 = cout_1931 ^ cout_1932; // @[Mul.scala 206:34]
  wire  cout_2029 = cout_1931 & cout_1932; // @[Mul.scala 207:34]
  wire  sum_2030 = sum_1935 ^ sum_1936; // @[Mul.scala 206:34]
  wire  cout_2030 = sum_1935 & sum_1936; // @[Mul.scala 207:34]
  wire  sum_2031 = cout_1933 ^ cout_1934; // @[Mul.scala 206:34]
  wire  cout_2031 = cout_1933 & cout_1934; // @[Mul.scala 207:34]
  wire  sum_2032 = sum_1937 ^ sum_1938; // @[Mul.scala 206:34]
  wire  cout_2032 = sum_1937 & sum_1938; // @[Mul.scala 207:34]
  wire  sum_2033 = cout_1935 ^ cout_1936; // @[Mul.scala 206:34]
  wire  cout_2033 = cout_1935 & cout_1936; // @[Mul.scala 207:34]
  wire  sum_2034 = sum_1939 ^ sum_1940; // @[Mul.scala 206:34]
  wire  cout_2034 = sum_1939 & sum_1940; // @[Mul.scala 207:34]
  wire  sum_2035 = cout_1937 ^ cout_1938; // @[Mul.scala 206:34]
  wire  cout_2035 = cout_1937 & cout_1938; // @[Mul.scala 207:34]
  wire  sum_2036 = sum_1941 ^ sum_1942; // @[Mul.scala 206:34]
  wire  cout_2036 = sum_1941 & sum_1942; // @[Mul.scala 207:34]
  wire  sum_2037 = cout_1939 ^ cout_1940; // @[Mul.scala 206:34]
  wire  cout_2037 = cout_1939 & cout_1940; // @[Mul.scala 207:34]
  wire  sum_2038 = sum_1943 ^ sum_1944; // @[Mul.scala 206:34]
  wire  cout_2038 = sum_1943 & sum_1944; // @[Mul.scala 207:34]
  wire  sum_2039 = cout_1941 ^ cout_1942; // @[Mul.scala 206:34]
  wire  cout_2039 = cout_1941 & cout_1942; // @[Mul.scala 207:34]
  wire  sum_2040 = sum_1945 ^ sum_1946; // @[Mul.scala 206:34]
  wire  cout_2040 = sum_1945 & sum_1946; // @[Mul.scala 207:34]
  wire  sum_2041 = cout_1943 ^ cout_1944; // @[Mul.scala 206:34]
  wire  cout_2041 = cout_1943 & cout_1944; // @[Mul.scala 207:34]
  wire  sum_2042 = sum_1947 ^ sum_1948; // @[Mul.scala 206:34]
  wire  cout_2042 = sum_1947 & sum_1948; // @[Mul.scala 207:34]
  wire  sum_2043 = cout_1945 ^ cout_1946; // @[Mul.scala 206:34]
  wire  cout_2043 = cout_1945 & cout_1946; // @[Mul.scala 207:34]
  wire  sum_2044 = sum_1949 ^ sum_1950; // @[Mul.scala 206:34]
  wire  cout_2044 = sum_1949 & sum_1950; // @[Mul.scala 207:34]
  wire  sum_2045 = cout_1947 ^ cout_1948; // @[Mul.scala 206:34]
  wire  cout_2045 = cout_1947 & cout_1948; // @[Mul.scala 207:34]
  wire  sum_2046 = sum_1951 ^ sum_1952; // @[Mul.scala 206:34]
  wire  cout_2046 = sum_1951 & sum_1952; // @[Mul.scala 207:34]
  wire  sum_2047 = cout_1949 ^ cout_1950; // @[Mul.scala 206:34]
  wire  cout_2047 = cout_1949 & cout_1950; // @[Mul.scala 207:34]
  wire  sum_2048 = sum_1953 ^ sum_1954; // @[Mul.scala 206:34]
  wire  cout_2048 = sum_1953 & sum_1954; // @[Mul.scala 207:34]
  wire  sum_2049 = cout_1951 ^ cout_1952; // @[Mul.scala 206:34]
  wire  cout_2049 = cout_1951 & cout_1952; // @[Mul.scala 207:34]
  wire  sum_2050 = sum_1955 ^ sum_1956; // @[Mul.scala 206:34]
  wire  cout_2050 = sum_1955 & sum_1956; // @[Mul.scala 207:34]
  wire  sum_2051 = cout_1953 ^ cout_1954; // @[Mul.scala 206:34]
  wire  cout_2051 = cout_1953 & cout_1954; // @[Mul.scala 207:34]
  wire  sum_2052 = sum_1957 ^ sum_1958; // @[Mul.scala 206:34]
  wire  cout_2052 = sum_1957 & sum_1958; // @[Mul.scala 207:34]
  wire  sum_2053 = cout_1955 ^ cout_1956; // @[Mul.scala 206:34]
  wire  cout_2053 = cout_1955 & cout_1956; // @[Mul.scala 207:34]
  wire  sum_2054 = sum_1959 ^ sum_1960; // @[Mul.scala 206:34]
  wire  cout_2054 = sum_1959 & sum_1960; // @[Mul.scala 207:34]
  wire  sum_2055 = cout_1957 ^ cout_1958; // @[Mul.scala 206:34]
  wire  cout_2055 = cout_1957 & cout_1958; // @[Mul.scala 207:34]
  wire  sum_2056 = sum_1961 ^ sum_1962; // @[Mul.scala 206:34]
  wire  cout_2056 = sum_1961 & sum_1962; // @[Mul.scala 207:34]
  wire  sum_2057 = cout_1959 ^ cout_1960; // @[Mul.scala 206:34]
  wire  cout_2057 = cout_1959 & cout_1960; // @[Mul.scala 207:34]
  wire  sum_2058 = sum_1963 ^ sum_1964; // @[Mul.scala 206:34]
  wire  cout_2058 = sum_1963 & sum_1964; // @[Mul.scala 207:34]
  wire  sum_2059 = cout_1961 ^ cout_1962; // @[Mul.scala 206:34]
  wire  cout_2059 = cout_1961 & cout_1962; // @[Mul.scala 207:34]
  wire  _sum_T_2700 = sum_1965 ^ cout_1963; // @[Mul.scala 191:34]
  wire  sum_2060 = sum_1965 ^ cout_1963 ^ cout_1964; // @[Mul.scala 191:42]
  wire  cout_2060 = sum_1965 & cout_1963 | _sum_T_2700 & cout_1964; // @[Mul.scala 192:44]
  wire  sum_2061 = sum_1966 ^ cout_1965; // @[Mul.scala 206:34]
  wire  cout_2061 = sum_1966 & cout_1965; // @[Mul.scala 207:34]
  wire  sum_2062 = sum_1967 ^ cout_1966; // @[Mul.scala 206:34]
  wire  cout_2062 = sum_1967 & cout_1966; // @[Mul.scala 207:34]
  wire  sum_2063 = sum_1968 ^ cout_1967; // @[Mul.scala 206:34]
  wire  cout_2063 = sum_1968 & cout_1967; // @[Mul.scala 207:34]
  wire  sum_2064 = sum_1969 ^ cout_1968; // @[Mul.scala 206:34]
  wire  cout_2064 = sum_1969 & cout_1968; // @[Mul.scala 207:34]
  wire  sum_2065 = sum_1970 ^ cout_1969; // @[Mul.scala 206:34]
  wire  sum_2088 = sum_1993 ^ cout_1992; // @[Mul.scala 206:34]
  wire  cout_2088 = sum_1993 & cout_1992; // @[Mul.scala 207:34]
  wire  sum_2089 = sum_1994 ^ cout_1993; // @[Mul.scala 206:34]
  wire  cout_2089 = sum_1994 & cout_1993; // @[Mul.scala 207:34]
  wire  sum_2090 = sum_1995 ^ cout_1994; // @[Mul.scala 206:34]
  wire  cout_2090 = sum_1995 & cout_1994; // @[Mul.scala 207:34]
  wire  _sum_T_2732 = sum_1996 ^ sum_1997; // @[Mul.scala 191:34]
  wire  sum_2091 = sum_1996 ^ sum_1997 ^ cout_1995; // @[Mul.scala 191:42]
  wire  cout_2091 = sum_1996 & sum_1997 | _sum_T_2732 & cout_1995; // @[Mul.scala 192:44]
  wire  sum_2092 = sum_1998 ^ sum_1999; // @[Mul.scala 206:34]
  wire  cout_2092 = sum_1998 & sum_1999; // @[Mul.scala 207:34]
  wire  sum_2093 = cout_1996 ^ cout_1997; // @[Mul.scala 206:34]
  wire  cout_2093 = cout_1996 & cout_1997; // @[Mul.scala 207:34]
  wire  sum_2094 = sum_2000 ^ sum_2001; // @[Mul.scala 206:34]
  wire  cout_2094 = sum_2000 & sum_2001; // @[Mul.scala 207:34]
  wire  sum_2095 = cout_1998 ^ cout_1999; // @[Mul.scala 206:34]
  wire  cout_2095 = cout_1998 & cout_1999; // @[Mul.scala 207:34]
  wire  sum_2096 = sum_2002 ^ sum_2003; // @[Mul.scala 206:34]
  wire  cout_2096 = sum_2002 & sum_2003; // @[Mul.scala 207:34]
  wire  sum_2097 = cout_2000 ^ cout_2001; // @[Mul.scala 206:34]
  wire  cout_2097 = cout_2000 & cout_2001; // @[Mul.scala 207:34]
  wire  sum_2098 = sum_2004 ^ sum_2005; // @[Mul.scala 206:34]
  wire  cout_2098 = sum_2004 & sum_2005; // @[Mul.scala 207:34]
  wire  sum_2099 = cout_2002 ^ cout_2003; // @[Mul.scala 206:34]
  wire  cout_2099 = cout_2002 & cout_2003; // @[Mul.scala 207:34]
  wire  sum_2100 = sum_2006 ^ sum_2007; // @[Mul.scala 206:34]
  wire  cout_2100 = sum_2006 & sum_2007; // @[Mul.scala 207:34]
  wire  sum_2101 = cout_2004 ^ cout_2005; // @[Mul.scala 206:34]
  wire  cout_2101 = cout_2004 & cout_2005; // @[Mul.scala 207:34]
  wire  sum_2102 = sum_2008 ^ sum_2009; // @[Mul.scala 206:34]
  wire  cout_2102 = sum_2008 & sum_2009; // @[Mul.scala 207:34]
  wire  sum_2103 = cout_2006 ^ cout_2007; // @[Mul.scala 206:34]
  wire  cout_2103 = cout_2006 & cout_2007; // @[Mul.scala 207:34]
  wire  sum_2104 = sum_2010 ^ sum_2011; // @[Mul.scala 206:34]
  wire  cout_2104 = sum_2010 & sum_2011; // @[Mul.scala 207:34]
  wire  sum_2105 = cout_2008 ^ cout_2009; // @[Mul.scala 206:34]
  wire  cout_2105 = cout_2008 & cout_2009; // @[Mul.scala 207:34]
  wire  sum_2106 = sum_2012 ^ sum_2013; // @[Mul.scala 206:34]
  wire  cout_2106 = sum_2012 & sum_2013; // @[Mul.scala 207:34]
  wire  sum_2107 = cout_2010 ^ cout_2011; // @[Mul.scala 206:34]
  wire  cout_2107 = cout_2010 & cout_2011; // @[Mul.scala 207:34]
  wire  sum_2108 = sum_2014 ^ sum_2015; // @[Mul.scala 206:34]
  wire  cout_2108 = sum_2014 & sum_2015; // @[Mul.scala 207:34]
  wire  sum_2109 = cout_2012 ^ cout_2013; // @[Mul.scala 206:34]
  wire  cout_2109 = cout_2012 & cout_2013; // @[Mul.scala 207:34]
  wire  sum_2110 = sum_2016 ^ sum_2017; // @[Mul.scala 206:34]
  wire  cout_2110 = sum_2016 & sum_2017; // @[Mul.scala 207:34]
  wire  sum_2111 = cout_2014 ^ cout_2015; // @[Mul.scala 206:34]
  wire  cout_2111 = cout_2014 & cout_2015; // @[Mul.scala 207:34]
  wire  sum_2112 = sum_2018 ^ sum_2019; // @[Mul.scala 206:34]
  wire  cout_2112 = sum_2018 & sum_2019; // @[Mul.scala 207:34]
  wire  sum_2113 = cout_2016 ^ cout_2017; // @[Mul.scala 206:34]
  wire  cout_2113 = cout_2016 & cout_2017; // @[Mul.scala 207:34]
  wire  sum_2114 = sum_2020 ^ sum_2021; // @[Mul.scala 206:34]
  wire  cout_2114 = sum_2020 & sum_2021; // @[Mul.scala 207:34]
  wire  sum_2115 = cout_2018 ^ cout_2019; // @[Mul.scala 206:34]
  wire  cout_2115 = cout_2018 & cout_2019; // @[Mul.scala 207:34]
  wire  sum_2116 = sum_2022 ^ sum_2023; // @[Mul.scala 206:34]
  wire  cout_2116 = sum_2022 & sum_2023; // @[Mul.scala 207:34]
  wire  sum_2117 = cout_2020 ^ cout_2021; // @[Mul.scala 206:34]
  wire  cout_2117 = cout_2020 & cout_2021; // @[Mul.scala 207:34]
  wire  sum_2118 = sum_2024 ^ sum_2025; // @[Mul.scala 206:34]
  wire  cout_2118 = sum_2024 & sum_2025; // @[Mul.scala 207:34]
  wire  sum_2119 = cout_2022 ^ cout_2023; // @[Mul.scala 206:34]
  wire  cout_2119 = cout_2022 & cout_2023; // @[Mul.scala 207:34]
  wire  sum_2120 = sum_2026 ^ sum_2027; // @[Mul.scala 206:34]
  wire  cout_2120 = sum_2026 & sum_2027; // @[Mul.scala 207:34]
  wire  sum_2121 = cout_2024 ^ cout_2025; // @[Mul.scala 206:34]
  wire  cout_2121 = cout_2024 & cout_2025; // @[Mul.scala 207:34]
  wire  sum_2122 = sum_2028 ^ sum_2029; // @[Mul.scala 206:34]
  wire  cout_2122 = sum_2028 & sum_2029; // @[Mul.scala 207:34]
  wire  sum_2123 = cout_2026 ^ cout_2027; // @[Mul.scala 206:34]
  wire  cout_2123 = cout_2026 & cout_2027; // @[Mul.scala 207:34]
  wire  sum_2124 = sum_2030 ^ sum_2031; // @[Mul.scala 206:34]
  wire  cout_2124 = sum_2030 & sum_2031; // @[Mul.scala 207:34]
  wire  sum_2125 = cout_2028 ^ cout_2029; // @[Mul.scala 206:34]
  wire  cout_2125 = cout_2028 & cout_2029; // @[Mul.scala 207:34]
  wire  sum_2126 = sum_2032 ^ sum_2033; // @[Mul.scala 206:34]
  wire  cout_2126 = sum_2032 & sum_2033; // @[Mul.scala 207:34]
  wire  sum_2127 = cout_2030 ^ cout_2031; // @[Mul.scala 206:34]
  wire  cout_2127 = cout_2030 & cout_2031; // @[Mul.scala 207:34]
  wire  sum_2128 = sum_2034 ^ sum_2035; // @[Mul.scala 206:34]
  wire  cout_2128 = sum_2034 & sum_2035; // @[Mul.scala 207:34]
  wire  sum_2129 = cout_2032 ^ cout_2033; // @[Mul.scala 206:34]
  wire  cout_2129 = cout_2032 & cout_2033; // @[Mul.scala 207:34]
  wire  sum_2130 = sum_2036 ^ sum_2037; // @[Mul.scala 206:34]
  wire  cout_2130 = sum_2036 & sum_2037; // @[Mul.scala 207:34]
  wire  sum_2131 = cout_2034 ^ cout_2035; // @[Mul.scala 206:34]
  wire  cout_2131 = cout_2034 & cout_2035; // @[Mul.scala 207:34]
  wire  sum_2132 = sum_2038 ^ sum_2039; // @[Mul.scala 206:34]
  wire  cout_2132 = sum_2038 & sum_2039; // @[Mul.scala 207:34]
  wire  sum_2133 = cout_2036 ^ cout_2037; // @[Mul.scala 206:34]
  wire  cout_2133 = cout_2036 & cout_2037; // @[Mul.scala 207:34]
  wire  sum_2134 = sum_2040 ^ sum_2041; // @[Mul.scala 206:34]
  wire  cout_2134 = sum_2040 & sum_2041; // @[Mul.scala 207:34]
  wire  sum_2135 = cout_2038 ^ cout_2039; // @[Mul.scala 206:34]
  wire  cout_2135 = cout_2038 & cout_2039; // @[Mul.scala 207:34]
  wire  sum_2136 = sum_2042 ^ sum_2043; // @[Mul.scala 206:34]
  wire  cout_2136 = sum_2042 & sum_2043; // @[Mul.scala 207:34]
  wire  sum_2137 = cout_2040 ^ cout_2041; // @[Mul.scala 206:34]
  wire  cout_2137 = cout_2040 & cout_2041; // @[Mul.scala 207:34]
  wire  sum_2138 = sum_2044 ^ sum_2045; // @[Mul.scala 206:34]
  wire  cout_2138 = sum_2044 & sum_2045; // @[Mul.scala 207:34]
  wire  sum_2139 = cout_2042 ^ cout_2043; // @[Mul.scala 206:34]
  wire  cout_2139 = cout_2042 & cout_2043; // @[Mul.scala 207:34]
  wire  sum_2140 = sum_2046 ^ sum_2047; // @[Mul.scala 206:34]
  wire  cout_2140 = sum_2046 & sum_2047; // @[Mul.scala 207:34]
  wire  sum_2141 = cout_2044 ^ cout_2045; // @[Mul.scala 206:34]
  wire  cout_2141 = cout_2044 & cout_2045; // @[Mul.scala 207:34]
  wire  sum_2142 = sum_2048 ^ sum_2049; // @[Mul.scala 206:34]
  wire  cout_2142 = sum_2048 & sum_2049; // @[Mul.scala 207:34]
  wire  sum_2143 = cout_2046 ^ cout_2047; // @[Mul.scala 206:34]
  wire  cout_2143 = cout_2046 & cout_2047; // @[Mul.scala 207:34]
  wire  sum_2144 = sum_2050 ^ sum_2051; // @[Mul.scala 206:34]
  wire  cout_2144 = sum_2050 & sum_2051; // @[Mul.scala 207:34]
  wire  sum_2145 = cout_2048 ^ cout_2049; // @[Mul.scala 206:34]
  wire  cout_2145 = cout_2048 & cout_2049; // @[Mul.scala 207:34]
  wire  sum_2146 = sum_2052 ^ sum_2053; // @[Mul.scala 206:34]
  wire  cout_2146 = sum_2052 & sum_2053; // @[Mul.scala 207:34]
  wire  sum_2147 = cout_2050 ^ cout_2051; // @[Mul.scala 206:34]
  wire  cout_2147 = cout_2050 & cout_2051; // @[Mul.scala 207:34]
  wire  sum_2148 = sum_2054 ^ sum_2055; // @[Mul.scala 206:34]
  wire  cout_2148 = sum_2054 & sum_2055; // @[Mul.scala 207:34]
  wire  sum_2149 = cout_2052 ^ cout_2053; // @[Mul.scala 206:34]
  wire  cout_2149 = cout_2052 & cout_2053; // @[Mul.scala 207:34]
  wire  sum_2150 = sum_2056 ^ sum_2057; // @[Mul.scala 206:34]
  wire  cout_2150 = sum_2056 & sum_2057; // @[Mul.scala 207:34]
  wire  sum_2151 = cout_2054 ^ cout_2055; // @[Mul.scala 206:34]
  wire  cout_2151 = cout_2054 & cout_2055; // @[Mul.scala 207:34]
  wire  sum_2152 = sum_2058 ^ sum_2059; // @[Mul.scala 206:34]
  wire  cout_2152 = sum_2058 & sum_2059; // @[Mul.scala 207:34]
  wire  sum_2153 = cout_2056 ^ cout_2057; // @[Mul.scala 206:34]
  wire  cout_2153 = cout_2056 & cout_2057; // @[Mul.scala 207:34]
  wire  _sum_T_2796 = sum_2060 ^ cout_2058; // @[Mul.scala 191:34]
  wire  sum_2154 = sum_2060 ^ cout_2058 ^ cout_2059; // @[Mul.scala 191:42]
  wire  cout_2154 = sum_2060 & cout_2058 | _sum_T_2796 & cout_2059; // @[Mul.scala 192:44]
  wire  sum_2155 = sum_2061 ^ cout_2060; // @[Mul.scala 206:34]
  wire  cout_2155 = sum_2061 & cout_2060; // @[Mul.scala 207:34]
  wire  sum_2156 = sum_2062 ^ cout_2061; // @[Mul.scala 206:34]
  wire  cout_2156 = sum_2062 & cout_2061; // @[Mul.scala 207:34]
  wire  sum_2157 = sum_2063 ^ cout_2062; // @[Mul.scala 206:34]
  wire  cout_2157 = sum_2063 & cout_2062; // @[Mul.scala 207:34]
  wire  sum_2158 = sum_2064 ^ cout_2063; // @[Mul.scala 206:34]
  wire  cout_2158 = sum_2064 & cout_2063; // @[Mul.scala 207:34]
  wire  sum_2159 = sum_2065 ^ cout_2064; // @[Mul.scala 206:34]
  wire  sum_2183 = sum_2089 ^ cout_2088; // @[Mul.scala 206:34]
  wire  cout_2183 = sum_2089 & cout_2088; // @[Mul.scala 207:34]
  wire  sum_2184 = sum_2090 ^ cout_2089; // @[Mul.scala 206:34]
  wire  cout_2184 = sum_2090 & cout_2089; // @[Mul.scala 207:34]
  wire  sum_2185 = sum_2091 ^ cout_2090; // @[Mul.scala 206:34]
  wire  cout_2185 = sum_2091 & cout_2090; // @[Mul.scala 207:34]
  wire  _sum_T_2829 = sum_2092 ^ sum_2093; // @[Mul.scala 191:34]
  wire  sum_2186 = sum_2092 ^ sum_2093 ^ cout_2091; // @[Mul.scala 191:42]
  wire  cout_2186 = sum_2092 & sum_2093 | _sum_T_2829 & cout_2091; // @[Mul.scala 192:44]
  wire  sum_2187 = sum_2094 ^ sum_2095; // @[Mul.scala 206:34]
  wire  cout_2187 = sum_2094 & sum_2095; // @[Mul.scala 207:34]
  wire  sum_2188 = cout_2092 ^ cout_2093; // @[Mul.scala 206:34]
  wire  cout_2188 = cout_2092 & cout_2093; // @[Mul.scala 207:34]
  wire  sum_2189 = sum_2096 ^ sum_2097; // @[Mul.scala 206:34]
  wire  cout_2189 = sum_2096 & sum_2097; // @[Mul.scala 207:34]
  wire  sum_2190 = cout_2094 ^ cout_2095; // @[Mul.scala 206:34]
  wire  cout_2190 = cout_2094 & cout_2095; // @[Mul.scala 207:34]
  wire  sum_2191 = sum_2098 ^ sum_2099; // @[Mul.scala 206:34]
  wire  cout_2191 = sum_2098 & sum_2099; // @[Mul.scala 207:34]
  wire  sum_2192 = cout_2096 ^ cout_2097; // @[Mul.scala 206:34]
  wire  cout_2192 = cout_2096 & cout_2097; // @[Mul.scala 207:34]
  wire  sum_2193 = sum_2100 ^ sum_2101; // @[Mul.scala 206:34]
  wire  cout_2193 = sum_2100 & sum_2101; // @[Mul.scala 207:34]
  wire  sum_2194 = cout_2098 ^ cout_2099; // @[Mul.scala 206:34]
  wire  cout_2194 = cout_2098 & cout_2099; // @[Mul.scala 207:34]
  wire  sum_2195 = sum_2102 ^ sum_2103; // @[Mul.scala 206:34]
  wire  cout_2195 = sum_2102 & sum_2103; // @[Mul.scala 207:34]
  wire  sum_2196 = cout_2100 ^ cout_2101; // @[Mul.scala 206:34]
  wire  cout_2196 = cout_2100 & cout_2101; // @[Mul.scala 207:34]
  wire  sum_2197 = sum_2104 ^ sum_2105; // @[Mul.scala 206:34]
  wire  cout_2197 = sum_2104 & sum_2105; // @[Mul.scala 207:34]
  wire  sum_2198 = cout_2102 ^ cout_2103; // @[Mul.scala 206:34]
  wire  cout_2198 = cout_2102 & cout_2103; // @[Mul.scala 207:34]
  wire  sum_2199 = sum_2106 ^ sum_2107; // @[Mul.scala 206:34]
  wire  cout_2199 = sum_2106 & sum_2107; // @[Mul.scala 207:34]
  wire  sum_2200 = cout_2104 ^ cout_2105; // @[Mul.scala 206:34]
  wire  cout_2200 = cout_2104 & cout_2105; // @[Mul.scala 207:34]
  wire  sum_2201 = sum_2108 ^ sum_2109; // @[Mul.scala 206:34]
  wire  cout_2201 = sum_2108 & sum_2109; // @[Mul.scala 207:34]
  wire  sum_2202 = cout_2106 ^ cout_2107; // @[Mul.scala 206:34]
  wire  cout_2202 = cout_2106 & cout_2107; // @[Mul.scala 207:34]
  wire  sum_2203 = sum_2110 ^ sum_2111; // @[Mul.scala 206:34]
  wire  cout_2203 = sum_2110 & sum_2111; // @[Mul.scala 207:34]
  wire  sum_2204 = cout_2108 ^ cout_2109; // @[Mul.scala 206:34]
  wire  cout_2204 = cout_2108 & cout_2109; // @[Mul.scala 207:34]
  wire  sum_2205 = sum_2112 ^ sum_2113; // @[Mul.scala 206:34]
  wire  cout_2205 = sum_2112 & sum_2113; // @[Mul.scala 207:34]
  wire  sum_2206 = cout_2110 ^ cout_2111; // @[Mul.scala 206:34]
  wire  cout_2206 = cout_2110 & cout_2111; // @[Mul.scala 207:34]
  wire  sum_2207 = sum_2114 ^ sum_2115; // @[Mul.scala 206:34]
  wire  cout_2207 = sum_2114 & sum_2115; // @[Mul.scala 207:34]
  wire  sum_2208 = cout_2112 ^ cout_2113; // @[Mul.scala 206:34]
  wire  cout_2208 = cout_2112 & cout_2113; // @[Mul.scala 207:34]
  wire  sum_2209 = sum_2116 ^ sum_2117; // @[Mul.scala 206:34]
  wire  cout_2209 = sum_2116 & sum_2117; // @[Mul.scala 207:34]
  wire  sum_2210 = cout_2114 ^ cout_2115; // @[Mul.scala 206:34]
  wire  cout_2210 = cout_2114 & cout_2115; // @[Mul.scala 207:34]
  wire  sum_2211 = sum_2118 ^ sum_2119; // @[Mul.scala 206:34]
  wire  cout_2211 = sum_2118 & sum_2119; // @[Mul.scala 207:34]
  wire  sum_2212 = cout_2116 ^ cout_2117; // @[Mul.scala 206:34]
  wire  cout_2212 = cout_2116 & cout_2117; // @[Mul.scala 207:34]
  wire  sum_2213 = sum_2120 ^ sum_2121; // @[Mul.scala 206:34]
  wire  cout_2213 = sum_2120 & sum_2121; // @[Mul.scala 207:34]
  wire  sum_2214 = cout_2118 ^ cout_2119; // @[Mul.scala 206:34]
  wire  cout_2214 = cout_2118 & cout_2119; // @[Mul.scala 207:34]
  wire  sum_2215 = sum_2122 ^ sum_2123; // @[Mul.scala 206:34]
  wire  cout_2215 = sum_2122 & sum_2123; // @[Mul.scala 207:34]
  wire  sum_2216 = cout_2120 ^ cout_2121; // @[Mul.scala 206:34]
  wire  cout_2216 = cout_2120 & cout_2121; // @[Mul.scala 207:34]
  wire  sum_2217 = sum_2124 ^ sum_2125; // @[Mul.scala 206:34]
  wire  cout_2217 = sum_2124 & sum_2125; // @[Mul.scala 207:34]
  wire  sum_2218 = cout_2122 ^ cout_2123; // @[Mul.scala 206:34]
  wire  cout_2218 = cout_2122 & cout_2123; // @[Mul.scala 207:34]
  wire  sum_2219 = sum_2126 ^ sum_2127; // @[Mul.scala 206:34]
  wire  cout_2219 = sum_2126 & sum_2127; // @[Mul.scala 207:34]
  wire  sum_2220 = cout_2124 ^ cout_2125; // @[Mul.scala 206:34]
  wire  cout_2220 = cout_2124 & cout_2125; // @[Mul.scala 207:34]
  wire  sum_2221 = sum_2128 ^ sum_2129; // @[Mul.scala 206:34]
  wire  cout_2221 = sum_2128 & sum_2129; // @[Mul.scala 207:34]
  wire  sum_2222 = cout_2126 ^ cout_2127; // @[Mul.scala 206:34]
  wire  cout_2222 = cout_2126 & cout_2127; // @[Mul.scala 207:34]
  wire  sum_2223 = sum_2130 ^ sum_2131; // @[Mul.scala 206:34]
  wire  cout_2223 = sum_2130 & sum_2131; // @[Mul.scala 207:34]
  wire  sum_2224 = cout_2128 ^ cout_2129; // @[Mul.scala 206:34]
  wire  cout_2224 = cout_2128 & cout_2129; // @[Mul.scala 207:34]
  wire  sum_2225 = sum_2132 ^ sum_2133; // @[Mul.scala 206:34]
  wire  cout_2225 = sum_2132 & sum_2133; // @[Mul.scala 207:34]
  wire  sum_2226 = cout_2130 ^ cout_2131; // @[Mul.scala 206:34]
  wire  cout_2226 = cout_2130 & cout_2131; // @[Mul.scala 207:34]
  wire  sum_2227 = sum_2134 ^ sum_2135; // @[Mul.scala 206:34]
  wire  cout_2227 = sum_2134 & sum_2135; // @[Mul.scala 207:34]
  wire  sum_2228 = cout_2132 ^ cout_2133; // @[Mul.scala 206:34]
  wire  cout_2228 = cout_2132 & cout_2133; // @[Mul.scala 207:34]
  wire  sum_2229 = sum_2136 ^ sum_2137; // @[Mul.scala 206:34]
  wire  cout_2229 = sum_2136 & sum_2137; // @[Mul.scala 207:34]
  wire  sum_2230 = cout_2134 ^ cout_2135; // @[Mul.scala 206:34]
  wire  cout_2230 = cout_2134 & cout_2135; // @[Mul.scala 207:34]
  wire  sum_2231 = sum_2138 ^ sum_2139; // @[Mul.scala 206:34]
  wire  cout_2231 = sum_2138 & sum_2139; // @[Mul.scala 207:34]
  wire  sum_2232 = cout_2136 ^ cout_2137; // @[Mul.scala 206:34]
  wire  cout_2232 = cout_2136 & cout_2137; // @[Mul.scala 207:34]
  wire  sum_2233 = sum_2140 ^ sum_2141; // @[Mul.scala 206:34]
  wire  cout_2233 = sum_2140 & sum_2141; // @[Mul.scala 207:34]
  wire  sum_2234 = cout_2138 ^ cout_2139; // @[Mul.scala 206:34]
  wire  cout_2234 = cout_2138 & cout_2139; // @[Mul.scala 207:34]
  wire  sum_2235 = sum_2142 ^ sum_2143; // @[Mul.scala 206:34]
  wire  cout_2235 = sum_2142 & sum_2143; // @[Mul.scala 207:34]
  wire  sum_2236 = cout_2140 ^ cout_2141; // @[Mul.scala 206:34]
  wire  cout_2236 = cout_2140 & cout_2141; // @[Mul.scala 207:34]
  wire  sum_2237 = sum_2144 ^ sum_2145; // @[Mul.scala 206:34]
  wire  cout_2237 = sum_2144 & sum_2145; // @[Mul.scala 207:34]
  wire  sum_2238 = cout_2142 ^ cout_2143; // @[Mul.scala 206:34]
  wire  cout_2238 = cout_2142 & cout_2143; // @[Mul.scala 207:34]
  wire  sum_2239 = sum_2146 ^ sum_2147; // @[Mul.scala 206:34]
  wire  cout_2239 = sum_2146 & sum_2147; // @[Mul.scala 207:34]
  wire  sum_2240 = cout_2144 ^ cout_2145; // @[Mul.scala 206:34]
  wire  cout_2240 = cout_2144 & cout_2145; // @[Mul.scala 207:34]
  wire  sum_2241 = sum_2148 ^ sum_2149; // @[Mul.scala 206:34]
  wire  cout_2241 = sum_2148 & sum_2149; // @[Mul.scala 207:34]
  wire  sum_2242 = cout_2146 ^ cout_2147; // @[Mul.scala 206:34]
  wire  cout_2242 = cout_2146 & cout_2147; // @[Mul.scala 207:34]
  wire  sum_2243 = sum_2150 ^ sum_2151; // @[Mul.scala 206:34]
  wire  cout_2243 = sum_2150 & sum_2151; // @[Mul.scala 207:34]
  wire  sum_2244 = cout_2148 ^ cout_2149; // @[Mul.scala 206:34]
  wire  cout_2244 = cout_2148 & cout_2149; // @[Mul.scala 207:34]
  wire  sum_2245 = sum_2152 ^ sum_2153; // @[Mul.scala 206:34]
  wire  cout_2245 = sum_2152 & sum_2153; // @[Mul.scala 207:34]
  wire  sum_2246 = cout_2150 ^ cout_2151; // @[Mul.scala 206:34]
  wire  cout_2246 = cout_2150 & cout_2151; // @[Mul.scala 207:34]
  wire  _sum_T_2891 = sum_2154 ^ cout_2152; // @[Mul.scala 191:34]
  wire  sum_2247 = sum_2154 ^ cout_2152 ^ cout_2153; // @[Mul.scala 191:42]
  wire  cout_2247 = sum_2154 & cout_2152 | _sum_T_2891 & cout_2153; // @[Mul.scala 192:44]
  wire  sum_2248 = sum_2155 ^ cout_2154; // @[Mul.scala 206:34]
  wire  cout_2248 = sum_2155 & cout_2154; // @[Mul.scala 207:34]
  wire  sum_2249 = sum_2156 ^ cout_2155; // @[Mul.scala 206:34]
  wire  cout_2249 = sum_2156 & cout_2155; // @[Mul.scala 207:34]
  wire  sum_2250 = sum_2157 ^ cout_2156; // @[Mul.scala 206:34]
  wire  cout_2250 = sum_2157 & cout_2156; // @[Mul.scala 207:34]
  wire  sum_2251 = sum_2158 ^ cout_2157; // @[Mul.scala 206:34]
  wire  cout_2251 = sum_2158 & cout_2157; // @[Mul.scala 207:34]
  wire  sum_2252 = sum_2159 ^ cout_2158; // @[Mul.scala 206:34]
  wire  sum_2277 = sum_2184 ^ cout_2183; // @[Mul.scala 206:34]
  wire  cout_2277 = sum_2184 & cout_2183; // @[Mul.scala 207:34]
  wire  sum_2278 = sum_2185 ^ cout_2184; // @[Mul.scala 206:34]
  wire  cout_2278 = sum_2185 & cout_2184; // @[Mul.scala 207:34]
  wire  sum_2279 = sum_2186 ^ cout_2185; // @[Mul.scala 206:34]
  wire  cout_2279 = sum_2186 & cout_2185; // @[Mul.scala 207:34]
  wire  _sum_T_2925 = sum_2187 ^ sum_2188; // @[Mul.scala 191:34]
  wire  sum_2280 = sum_2187 ^ sum_2188 ^ cout_2186; // @[Mul.scala 191:42]
  wire  cout_2280 = sum_2187 & sum_2188 | _sum_T_2925 & cout_2186; // @[Mul.scala 192:44]
  wire  sum_2281 = sum_2189 ^ sum_2190; // @[Mul.scala 206:34]
  wire  cout_2281 = sum_2189 & sum_2190; // @[Mul.scala 207:34]
  wire  sum_2282 = cout_2187 ^ cout_2188; // @[Mul.scala 206:34]
  wire  cout_2282 = cout_2187 & cout_2188; // @[Mul.scala 207:34]
  wire  sum_2283 = sum_2191 ^ sum_2192; // @[Mul.scala 206:34]
  wire  cout_2283 = sum_2191 & sum_2192; // @[Mul.scala 207:34]
  wire  sum_2284 = cout_2189 ^ cout_2190; // @[Mul.scala 206:34]
  wire  cout_2284 = cout_2189 & cout_2190; // @[Mul.scala 207:34]
  wire  sum_2285 = sum_2193 ^ sum_2194; // @[Mul.scala 206:34]
  wire  cout_2285 = sum_2193 & sum_2194; // @[Mul.scala 207:34]
  wire  sum_2286 = cout_2191 ^ cout_2192; // @[Mul.scala 206:34]
  wire  cout_2286 = cout_2191 & cout_2192; // @[Mul.scala 207:34]
  wire  sum_2287 = sum_2195 ^ sum_2196; // @[Mul.scala 206:34]
  wire  cout_2287 = sum_2195 & sum_2196; // @[Mul.scala 207:34]
  wire  sum_2288 = cout_2193 ^ cout_2194; // @[Mul.scala 206:34]
  wire  cout_2288 = cout_2193 & cout_2194; // @[Mul.scala 207:34]
  wire  sum_2289 = sum_2197 ^ sum_2198; // @[Mul.scala 206:34]
  wire  cout_2289 = sum_2197 & sum_2198; // @[Mul.scala 207:34]
  wire  sum_2290 = cout_2195 ^ cout_2196; // @[Mul.scala 206:34]
  wire  cout_2290 = cout_2195 & cout_2196; // @[Mul.scala 207:34]
  wire  sum_2291 = sum_2199 ^ sum_2200; // @[Mul.scala 206:34]
  wire  cout_2291 = sum_2199 & sum_2200; // @[Mul.scala 207:34]
  wire  sum_2292 = cout_2197 ^ cout_2198; // @[Mul.scala 206:34]
  wire  cout_2292 = cout_2197 & cout_2198; // @[Mul.scala 207:34]
  wire  sum_2293 = sum_2201 ^ sum_2202; // @[Mul.scala 206:34]
  wire  cout_2293 = sum_2201 & sum_2202; // @[Mul.scala 207:34]
  wire  sum_2294 = cout_2199 ^ cout_2200; // @[Mul.scala 206:34]
  wire  cout_2294 = cout_2199 & cout_2200; // @[Mul.scala 207:34]
  wire  sum_2295 = sum_2203 ^ sum_2204; // @[Mul.scala 206:34]
  wire  cout_2295 = sum_2203 & sum_2204; // @[Mul.scala 207:34]
  wire  sum_2296 = cout_2201 ^ cout_2202; // @[Mul.scala 206:34]
  wire  cout_2296 = cout_2201 & cout_2202; // @[Mul.scala 207:34]
  wire  sum_2297 = sum_2205 ^ sum_2206; // @[Mul.scala 206:34]
  wire  cout_2297 = sum_2205 & sum_2206; // @[Mul.scala 207:34]
  wire  sum_2298 = cout_2203 ^ cout_2204; // @[Mul.scala 206:34]
  wire  cout_2298 = cout_2203 & cout_2204; // @[Mul.scala 207:34]
  wire  sum_2299 = sum_2207 ^ sum_2208; // @[Mul.scala 206:34]
  wire  cout_2299 = sum_2207 & sum_2208; // @[Mul.scala 207:34]
  wire  sum_2300 = cout_2205 ^ cout_2206; // @[Mul.scala 206:34]
  wire  cout_2300 = cout_2205 & cout_2206; // @[Mul.scala 207:34]
  wire  sum_2301 = sum_2209 ^ sum_2210; // @[Mul.scala 206:34]
  wire  cout_2301 = sum_2209 & sum_2210; // @[Mul.scala 207:34]
  wire  sum_2302 = cout_2207 ^ cout_2208; // @[Mul.scala 206:34]
  wire  cout_2302 = cout_2207 & cout_2208; // @[Mul.scala 207:34]
  wire  sum_2303 = sum_2211 ^ sum_2212; // @[Mul.scala 206:34]
  wire  cout_2303 = sum_2211 & sum_2212; // @[Mul.scala 207:34]
  wire  sum_2304 = cout_2209 ^ cout_2210; // @[Mul.scala 206:34]
  wire  cout_2304 = cout_2209 & cout_2210; // @[Mul.scala 207:34]
  wire  sum_2305 = sum_2213 ^ sum_2214; // @[Mul.scala 206:34]
  wire  cout_2305 = sum_2213 & sum_2214; // @[Mul.scala 207:34]
  wire  sum_2306 = cout_2211 ^ cout_2212; // @[Mul.scala 206:34]
  wire  cout_2306 = cout_2211 & cout_2212; // @[Mul.scala 207:34]
  wire  sum_2307 = sum_2215 ^ sum_2216; // @[Mul.scala 206:34]
  wire  cout_2307 = sum_2215 & sum_2216; // @[Mul.scala 207:34]
  wire  sum_2308 = cout_2213 ^ cout_2214; // @[Mul.scala 206:34]
  wire  cout_2308 = cout_2213 & cout_2214; // @[Mul.scala 207:34]
  wire  sum_2309 = sum_2217 ^ sum_2218; // @[Mul.scala 206:34]
  wire  cout_2309 = sum_2217 & sum_2218; // @[Mul.scala 207:34]
  wire  sum_2310 = cout_2215 ^ cout_2216; // @[Mul.scala 206:34]
  wire  cout_2310 = cout_2215 & cout_2216; // @[Mul.scala 207:34]
  wire  sum_2311 = sum_2219 ^ sum_2220; // @[Mul.scala 206:34]
  wire  cout_2311 = sum_2219 & sum_2220; // @[Mul.scala 207:34]
  wire  sum_2312 = cout_2217 ^ cout_2218; // @[Mul.scala 206:34]
  wire  cout_2312 = cout_2217 & cout_2218; // @[Mul.scala 207:34]
  wire  sum_2313 = sum_2221 ^ sum_2222; // @[Mul.scala 206:34]
  wire  cout_2313 = sum_2221 & sum_2222; // @[Mul.scala 207:34]
  wire  sum_2314 = cout_2219 ^ cout_2220; // @[Mul.scala 206:34]
  wire  cout_2314 = cout_2219 & cout_2220; // @[Mul.scala 207:34]
  wire  sum_2315 = sum_2223 ^ sum_2224; // @[Mul.scala 206:34]
  wire  cout_2315 = sum_2223 & sum_2224; // @[Mul.scala 207:34]
  wire  sum_2316 = cout_2221 ^ cout_2222; // @[Mul.scala 206:34]
  wire  cout_2316 = cout_2221 & cout_2222; // @[Mul.scala 207:34]
  wire  sum_2317 = sum_2225 ^ sum_2226; // @[Mul.scala 206:34]
  wire  cout_2317 = sum_2225 & sum_2226; // @[Mul.scala 207:34]
  wire  sum_2318 = cout_2223 ^ cout_2224; // @[Mul.scala 206:34]
  wire  cout_2318 = cout_2223 & cout_2224; // @[Mul.scala 207:34]
  wire  sum_2319 = sum_2227 ^ sum_2228; // @[Mul.scala 206:34]
  wire  cout_2319 = sum_2227 & sum_2228; // @[Mul.scala 207:34]
  wire  sum_2320 = cout_2225 ^ cout_2226; // @[Mul.scala 206:34]
  wire  cout_2320 = cout_2225 & cout_2226; // @[Mul.scala 207:34]
  wire  sum_2321 = sum_2229 ^ sum_2230; // @[Mul.scala 206:34]
  wire  cout_2321 = sum_2229 & sum_2230; // @[Mul.scala 207:34]
  wire  sum_2322 = cout_2227 ^ cout_2228; // @[Mul.scala 206:34]
  wire  cout_2322 = cout_2227 & cout_2228; // @[Mul.scala 207:34]
  wire  sum_2323 = sum_2231 ^ sum_2232; // @[Mul.scala 206:34]
  wire  cout_2323 = sum_2231 & sum_2232; // @[Mul.scala 207:34]
  wire  sum_2324 = cout_2229 ^ cout_2230; // @[Mul.scala 206:34]
  wire  cout_2324 = cout_2229 & cout_2230; // @[Mul.scala 207:34]
  wire  sum_2325 = sum_2233 ^ sum_2234; // @[Mul.scala 206:34]
  wire  cout_2325 = sum_2233 & sum_2234; // @[Mul.scala 207:34]
  wire  sum_2326 = cout_2231 ^ cout_2232; // @[Mul.scala 206:34]
  wire  cout_2326 = cout_2231 & cout_2232; // @[Mul.scala 207:34]
  wire  sum_2327 = sum_2235 ^ sum_2236; // @[Mul.scala 206:34]
  wire  cout_2327 = sum_2235 & sum_2236; // @[Mul.scala 207:34]
  wire  sum_2328 = cout_2233 ^ cout_2234; // @[Mul.scala 206:34]
  wire  cout_2328 = cout_2233 & cout_2234; // @[Mul.scala 207:34]
  wire  sum_2329 = sum_2237 ^ sum_2238; // @[Mul.scala 206:34]
  wire  cout_2329 = sum_2237 & sum_2238; // @[Mul.scala 207:34]
  wire  sum_2330 = cout_2235 ^ cout_2236; // @[Mul.scala 206:34]
  wire  cout_2330 = cout_2235 & cout_2236; // @[Mul.scala 207:34]
  wire  sum_2331 = sum_2239 ^ sum_2240; // @[Mul.scala 206:34]
  wire  cout_2331 = sum_2239 & sum_2240; // @[Mul.scala 207:34]
  wire  sum_2332 = cout_2237 ^ cout_2238; // @[Mul.scala 206:34]
  wire  cout_2332 = cout_2237 & cout_2238; // @[Mul.scala 207:34]
  wire  sum_2333 = sum_2241 ^ sum_2242; // @[Mul.scala 206:34]
  wire  cout_2333 = sum_2241 & sum_2242; // @[Mul.scala 207:34]
  wire  sum_2334 = cout_2239 ^ cout_2240; // @[Mul.scala 206:34]
  wire  cout_2334 = cout_2239 & cout_2240; // @[Mul.scala 207:34]
  wire  sum_2335 = sum_2243 ^ sum_2244; // @[Mul.scala 206:34]
  wire  cout_2335 = sum_2243 & sum_2244; // @[Mul.scala 207:34]
  wire  sum_2336 = cout_2241 ^ cout_2242; // @[Mul.scala 206:34]
  wire  cout_2336 = cout_2241 & cout_2242; // @[Mul.scala 207:34]
  wire  sum_2337 = sum_2245 ^ sum_2246; // @[Mul.scala 206:34]
  wire  cout_2337 = sum_2245 & sum_2246; // @[Mul.scala 207:34]
  wire  sum_2338 = cout_2243 ^ cout_2244; // @[Mul.scala 206:34]
  wire  cout_2338 = cout_2243 & cout_2244; // @[Mul.scala 207:34]
  wire  _sum_T_2985 = sum_2247 ^ cout_2245; // @[Mul.scala 191:34]
  wire  sum_2339 = sum_2247 ^ cout_2245 ^ cout_2246; // @[Mul.scala 191:42]
  wire  cout_2339 = sum_2247 & cout_2245 | _sum_T_2985 & cout_2246; // @[Mul.scala 192:44]
  wire  sum_2340 = sum_2248 ^ cout_2247; // @[Mul.scala 206:34]
  wire  cout_2340 = sum_2248 & cout_2247; // @[Mul.scala 207:34]
  wire  sum_2341 = sum_2249 ^ cout_2248; // @[Mul.scala 206:34]
  wire  cout_2341 = sum_2249 & cout_2248; // @[Mul.scala 207:34]
  wire  sum_2342 = sum_2250 ^ cout_2249; // @[Mul.scala 206:34]
  wire  cout_2342 = sum_2250 & cout_2249; // @[Mul.scala 207:34]
  wire  sum_2343 = sum_2251 ^ cout_2250; // @[Mul.scala 206:34]
  wire  cout_2343 = sum_2251 & cout_2250; // @[Mul.scala 207:34]
  wire  sum_2344 = sum_2252 ^ cout_2251; // @[Mul.scala 206:34]
  wire  sum_2370 = sum_2278 ^ cout_2277; // @[Mul.scala 206:34]
  wire  cout_2370 = sum_2278 & cout_2277; // @[Mul.scala 207:34]
  wire  sum_2371 = sum_2279 ^ cout_2278; // @[Mul.scala 206:34]
  wire  cout_2371 = sum_2279 & cout_2278; // @[Mul.scala 207:34]
  wire  sum_2372 = sum_2280 ^ cout_2279; // @[Mul.scala 206:34]
  wire  cout_2372 = sum_2280 & cout_2279; // @[Mul.scala 207:34]
  wire  _sum_T_3020 = sum_2281 ^ sum_2282; // @[Mul.scala 191:34]
  wire  sum_2373 = sum_2281 ^ sum_2282 ^ cout_2280; // @[Mul.scala 191:42]
  wire  cout_2373 = sum_2281 & sum_2282 | _sum_T_3020 & cout_2280; // @[Mul.scala 192:44]
  wire  sum_2374 = sum_2283 ^ sum_2284; // @[Mul.scala 206:34]
  wire  cout_2374 = sum_2283 & sum_2284; // @[Mul.scala 207:34]
  wire  sum_2375 = cout_2281 ^ cout_2282; // @[Mul.scala 206:34]
  wire  cout_2375 = cout_2281 & cout_2282; // @[Mul.scala 207:34]
  wire  sum_2376 = sum_2285 ^ sum_2286; // @[Mul.scala 206:34]
  wire  cout_2376 = sum_2285 & sum_2286; // @[Mul.scala 207:34]
  wire  sum_2377 = cout_2283 ^ cout_2284; // @[Mul.scala 206:34]
  wire  cout_2377 = cout_2283 & cout_2284; // @[Mul.scala 207:34]
  wire  sum_2378 = sum_2287 ^ sum_2288; // @[Mul.scala 206:34]
  wire  cout_2378 = sum_2287 & sum_2288; // @[Mul.scala 207:34]
  wire  sum_2379 = cout_2285 ^ cout_2286; // @[Mul.scala 206:34]
  wire  cout_2379 = cout_2285 & cout_2286; // @[Mul.scala 207:34]
  wire  sum_2380 = sum_2289 ^ sum_2290; // @[Mul.scala 206:34]
  wire  cout_2380 = sum_2289 & sum_2290; // @[Mul.scala 207:34]
  wire  sum_2381 = cout_2287 ^ cout_2288; // @[Mul.scala 206:34]
  wire  cout_2381 = cout_2287 & cout_2288; // @[Mul.scala 207:34]
  wire  sum_2382 = sum_2291 ^ sum_2292; // @[Mul.scala 206:34]
  wire  cout_2382 = sum_2291 & sum_2292; // @[Mul.scala 207:34]
  wire  sum_2383 = cout_2289 ^ cout_2290; // @[Mul.scala 206:34]
  wire  cout_2383 = cout_2289 & cout_2290; // @[Mul.scala 207:34]
  wire  sum_2384 = sum_2293 ^ sum_2294; // @[Mul.scala 206:34]
  wire  cout_2384 = sum_2293 & sum_2294; // @[Mul.scala 207:34]
  wire  sum_2385 = cout_2291 ^ cout_2292; // @[Mul.scala 206:34]
  wire  cout_2385 = cout_2291 & cout_2292; // @[Mul.scala 207:34]
  wire  sum_2386 = sum_2295 ^ sum_2296; // @[Mul.scala 206:34]
  wire  cout_2386 = sum_2295 & sum_2296; // @[Mul.scala 207:34]
  wire  sum_2387 = cout_2293 ^ cout_2294; // @[Mul.scala 206:34]
  wire  cout_2387 = cout_2293 & cout_2294; // @[Mul.scala 207:34]
  wire  sum_2388 = sum_2297 ^ sum_2298; // @[Mul.scala 206:34]
  wire  cout_2388 = sum_2297 & sum_2298; // @[Mul.scala 207:34]
  wire  sum_2389 = cout_2295 ^ cout_2296; // @[Mul.scala 206:34]
  wire  cout_2389 = cout_2295 & cout_2296; // @[Mul.scala 207:34]
  wire  sum_2390 = sum_2299 ^ sum_2300; // @[Mul.scala 206:34]
  wire  cout_2390 = sum_2299 & sum_2300; // @[Mul.scala 207:34]
  wire  sum_2391 = cout_2297 ^ cout_2298; // @[Mul.scala 206:34]
  wire  cout_2391 = cout_2297 & cout_2298; // @[Mul.scala 207:34]
  wire  sum_2392 = sum_2301 ^ sum_2302; // @[Mul.scala 206:34]
  wire  cout_2392 = sum_2301 & sum_2302; // @[Mul.scala 207:34]
  wire  sum_2393 = cout_2299 ^ cout_2300; // @[Mul.scala 206:34]
  wire  cout_2393 = cout_2299 & cout_2300; // @[Mul.scala 207:34]
  wire  sum_2394 = sum_2303 ^ sum_2304; // @[Mul.scala 206:34]
  wire  cout_2394 = sum_2303 & sum_2304; // @[Mul.scala 207:34]
  wire  sum_2395 = cout_2301 ^ cout_2302; // @[Mul.scala 206:34]
  wire  cout_2395 = cout_2301 & cout_2302; // @[Mul.scala 207:34]
  wire  sum_2396 = sum_2305 ^ sum_2306; // @[Mul.scala 206:34]
  wire  cout_2396 = sum_2305 & sum_2306; // @[Mul.scala 207:34]
  wire  sum_2397 = cout_2303 ^ cout_2304; // @[Mul.scala 206:34]
  wire  cout_2397 = cout_2303 & cout_2304; // @[Mul.scala 207:34]
  wire  sum_2398 = sum_2307 ^ sum_2308; // @[Mul.scala 206:34]
  wire  cout_2398 = sum_2307 & sum_2308; // @[Mul.scala 207:34]
  wire  sum_2399 = cout_2305 ^ cout_2306; // @[Mul.scala 206:34]
  wire  cout_2399 = cout_2305 & cout_2306; // @[Mul.scala 207:34]
  wire  sum_2400 = sum_2309 ^ sum_2310; // @[Mul.scala 206:34]
  wire  cout_2400 = sum_2309 & sum_2310; // @[Mul.scala 207:34]
  wire  sum_2401 = cout_2307 ^ cout_2308; // @[Mul.scala 206:34]
  wire  cout_2401 = cout_2307 & cout_2308; // @[Mul.scala 207:34]
  wire  sum_2402 = sum_2311 ^ sum_2312; // @[Mul.scala 206:34]
  wire  cout_2402 = sum_2311 & sum_2312; // @[Mul.scala 207:34]
  wire  sum_2403 = cout_2309 ^ cout_2310; // @[Mul.scala 206:34]
  wire  cout_2403 = cout_2309 & cout_2310; // @[Mul.scala 207:34]
  wire  sum_2404 = sum_2313 ^ sum_2314; // @[Mul.scala 206:34]
  wire  cout_2404 = sum_2313 & sum_2314; // @[Mul.scala 207:34]
  wire  sum_2405 = cout_2311 ^ cout_2312; // @[Mul.scala 206:34]
  wire  cout_2405 = cout_2311 & cout_2312; // @[Mul.scala 207:34]
  wire  sum_2406 = sum_2315 ^ sum_2316; // @[Mul.scala 206:34]
  wire  cout_2406 = sum_2315 & sum_2316; // @[Mul.scala 207:34]
  wire  sum_2407 = cout_2313 ^ cout_2314; // @[Mul.scala 206:34]
  wire  cout_2407 = cout_2313 & cout_2314; // @[Mul.scala 207:34]
  wire  sum_2408 = sum_2317 ^ sum_2318; // @[Mul.scala 206:34]
  wire  cout_2408 = sum_2317 & sum_2318; // @[Mul.scala 207:34]
  wire  sum_2409 = cout_2315 ^ cout_2316; // @[Mul.scala 206:34]
  wire  cout_2409 = cout_2315 & cout_2316; // @[Mul.scala 207:34]
  wire  sum_2410 = sum_2319 ^ sum_2320; // @[Mul.scala 206:34]
  wire  cout_2410 = sum_2319 & sum_2320; // @[Mul.scala 207:34]
  wire  sum_2411 = cout_2317 ^ cout_2318; // @[Mul.scala 206:34]
  wire  cout_2411 = cout_2317 & cout_2318; // @[Mul.scala 207:34]
  wire  sum_2412 = sum_2321 ^ sum_2322; // @[Mul.scala 206:34]
  wire  cout_2412 = sum_2321 & sum_2322; // @[Mul.scala 207:34]
  wire  sum_2413 = cout_2319 ^ cout_2320; // @[Mul.scala 206:34]
  wire  cout_2413 = cout_2319 & cout_2320; // @[Mul.scala 207:34]
  wire  sum_2414 = sum_2323 ^ sum_2324; // @[Mul.scala 206:34]
  wire  cout_2414 = sum_2323 & sum_2324; // @[Mul.scala 207:34]
  wire  sum_2415 = cout_2321 ^ cout_2322; // @[Mul.scala 206:34]
  wire  cout_2415 = cout_2321 & cout_2322; // @[Mul.scala 207:34]
  wire  sum_2416 = sum_2325 ^ sum_2326; // @[Mul.scala 206:34]
  wire  cout_2416 = sum_2325 & sum_2326; // @[Mul.scala 207:34]
  wire  sum_2417 = cout_2323 ^ cout_2324; // @[Mul.scala 206:34]
  wire  cout_2417 = cout_2323 & cout_2324; // @[Mul.scala 207:34]
  wire  sum_2418 = sum_2327 ^ sum_2328; // @[Mul.scala 206:34]
  wire  cout_2418 = sum_2327 & sum_2328; // @[Mul.scala 207:34]
  wire  sum_2419 = cout_2325 ^ cout_2326; // @[Mul.scala 206:34]
  wire  cout_2419 = cout_2325 & cout_2326; // @[Mul.scala 207:34]
  wire  sum_2420 = sum_2329 ^ sum_2330; // @[Mul.scala 206:34]
  wire  cout_2420 = sum_2329 & sum_2330; // @[Mul.scala 207:34]
  wire  sum_2421 = cout_2327 ^ cout_2328; // @[Mul.scala 206:34]
  wire  cout_2421 = cout_2327 & cout_2328; // @[Mul.scala 207:34]
  wire  sum_2422 = sum_2331 ^ sum_2332; // @[Mul.scala 206:34]
  wire  cout_2422 = sum_2331 & sum_2332; // @[Mul.scala 207:34]
  wire  sum_2423 = cout_2329 ^ cout_2330; // @[Mul.scala 206:34]
  wire  cout_2423 = cout_2329 & cout_2330; // @[Mul.scala 207:34]
  wire  sum_2424 = sum_2333 ^ sum_2334; // @[Mul.scala 206:34]
  wire  cout_2424 = sum_2333 & sum_2334; // @[Mul.scala 207:34]
  wire  sum_2425 = cout_2331 ^ cout_2332; // @[Mul.scala 206:34]
  wire  cout_2425 = cout_2331 & cout_2332; // @[Mul.scala 207:34]
  wire  sum_2426 = sum_2335 ^ sum_2336; // @[Mul.scala 206:34]
  wire  cout_2426 = sum_2335 & sum_2336; // @[Mul.scala 207:34]
  wire  sum_2427 = cout_2333 ^ cout_2334; // @[Mul.scala 206:34]
  wire  cout_2427 = cout_2333 & cout_2334; // @[Mul.scala 207:34]
  wire  sum_2428 = sum_2337 ^ sum_2338; // @[Mul.scala 206:34]
  wire  cout_2428 = sum_2337 & sum_2338; // @[Mul.scala 207:34]
  wire  sum_2429 = cout_2335 ^ cout_2336; // @[Mul.scala 206:34]
  wire  cout_2429 = cout_2335 & cout_2336; // @[Mul.scala 207:34]
  wire  _sum_T_3078 = sum_2339 ^ cout_2337; // @[Mul.scala 191:34]
  wire  sum_2430 = sum_2339 ^ cout_2337 ^ cout_2338; // @[Mul.scala 191:42]
  wire  cout_2430 = sum_2339 & cout_2337 | _sum_T_3078 & cout_2338; // @[Mul.scala 192:44]
  wire  sum_2431 = sum_2340 ^ cout_2339; // @[Mul.scala 206:34]
  wire  cout_2431 = sum_2340 & cout_2339; // @[Mul.scala 207:34]
  wire  sum_2432 = sum_2341 ^ cout_2340; // @[Mul.scala 206:34]
  wire  cout_2432 = sum_2341 & cout_2340; // @[Mul.scala 207:34]
  wire  sum_2433 = sum_2342 ^ cout_2341; // @[Mul.scala 206:34]
  wire  cout_2433 = sum_2342 & cout_2341; // @[Mul.scala 207:34]
  wire  sum_2434 = sum_2343 ^ cout_2342; // @[Mul.scala 206:34]
  wire  cout_2434 = sum_2343 & cout_2342; // @[Mul.scala 207:34]
  wire  sum_2435 = sum_2344 ^ cout_2343; // @[Mul.scala 206:34]
  wire  sum_2462 = sum_2371 ^ cout_2370; // @[Mul.scala 206:34]
  wire  cout_2462 = sum_2371 & cout_2370; // @[Mul.scala 207:34]
  wire  sum_2463 = sum_2372 ^ cout_2371; // @[Mul.scala 206:34]
  wire  cout_2463 = sum_2372 & cout_2371; // @[Mul.scala 207:34]
  wire  sum_2464 = sum_2373 ^ cout_2372; // @[Mul.scala 206:34]
  wire  cout_2464 = sum_2373 & cout_2372; // @[Mul.scala 207:34]
  wire  _sum_T_3114 = sum_2374 ^ sum_2375; // @[Mul.scala 191:34]
  wire  sum_2465 = sum_2374 ^ sum_2375 ^ cout_2373; // @[Mul.scala 191:42]
  wire  cout_2465 = sum_2374 & sum_2375 | _sum_T_3114 & cout_2373; // @[Mul.scala 192:44]
  wire  sum_2466 = sum_2376 ^ sum_2377; // @[Mul.scala 206:34]
  wire  cout_2466 = sum_2376 & sum_2377; // @[Mul.scala 207:34]
  wire  sum_2467 = cout_2374 ^ cout_2375; // @[Mul.scala 206:34]
  wire  cout_2467 = cout_2374 & cout_2375; // @[Mul.scala 207:34]
  wire  sum_2468 = sum_2378 ^ sum_2379; // @[Mul.scala 206:34]
  wire  cout_2468 = sum_2378 & sum_2379; // @[Mul.scala 207:34]
  wire  sum_2469 = cout_2376 ^ cout_2377; // @[Mul.scala 206:34]
  wire  cout_2469 = cout_2376 & cout_2377; // @[Mul.scala 207:34]
  wire  sum_2470 = sum_2380 ^ sum_2381; // @[Mul.scala 206:34]
  wire  cout_2470 = sum_2380 & sum_2381; // @[Mul.scala 207:34]
  wire  sum_2471 = cout_2378 ^ cout_2379; // @[Mul.scala 206:34]
  wire  cout_2471 = cout_2378 & cout_2379; // @[Mul.scala 207:34]
  wire  sum_2472 = sum_2382 ^ sum_2383; // @[Mul.scala 206:34]
  wire  cout_2472 = sum_2382 & sum_2383; // @[Mul.scala 207:34]
  wire  sum_2473 = cout_2380 ^ cout_2381; // @[Mul.scala 206:34]
  wire  cout_2473 = cout_2380 & cout_2381; // @[Mul.scala 207:34]
  wire  sum_2474 = sum_2384 ^ sum_2385; // @[Mul.scala 206:34]
  wire  cout_2474 = sum_2384 & sum_2385; // @[Mul.scala 207:34]
  wire  sum_2475 = cout_2382 ^ cout_2383; // @[Mul.scala 206:34]
  wire  cout_2475 = cout_2382 & cout_2383; // @[Mul.scala 207:34]
  wire  sum_2476 = sum_2386 ^ sum_2387; // @[Mul.scala 206:34]
  wire  cout_2476 = sum_2386 & sum_2387; // @[Mul.scala 207:34]
  wire  sum_2477 = cout_2384 ^ cout_2385; // @[Mul.scala 206:34]
  wire  cout_2477 = cout_2384 & cout_2385; // @[Mul.scala 207:34]
  wire  sum_2478 = sum_2388 ^ sum_2389; // @[Mul.scala 206:34]
  wire  cout_2478 = sum_2388 & sum_2389; // @[Mul.scala 207:34]
  wire  sum_2479 = cout_2386 ^ cout_2387; // @[Mul.scala 206:34]
  wire  cout_2479 = cout_2386 & cout_2387; // @[Mul.scala 207:34]
  wire  sum_2480 = sum_2390 ^ sum_2391; // @[Mul.scala 206:34]
  wire  cout_2480 = sum_2390 & sum_2391; // @[Mul.scala 207:34]
  wire  sum_2481 = cout_2388 ^ cout_2389; // @[Mul.scala 206:34]
  wire  cout_2481 = cout_2388 & cout_2389; // @[Mul.scala 207:34]
  wire  sum_2482 = sum_2392 ^ sum_2393; // @[Mul.scala 206:34]
  wire  cout_2482 = sum_2392 & sum_2393; // @[Mul.scala 207:34]
  wire  sum_2483 = cout_2390 ^ cout_2391; // @[Mul.scala 206:34]
  wire  cout_2483 = cout_2390 & cout_2391; // @[Mul.scala 207:34]
  wire  sum_2484 = sum_2394 ^ sum_2395; // @[Mul.scala 206:34]
  wire  cout_2484 = sum_2394 & sum_2395; // @[Mul.scala 207:34]
  wire  sum_2485 = cout_2392 ^ cout_2393; // @[Mul.scala 206:34]
  wire  cout_2485 = cout_2392 & cout_2393; // @[Mul.scala 207:34]
  wire  sum_2486 = sum_2396 ^ sum_2397; // @[Mul.scala 206:34]
  wire  cout_2486 = sum_2396 & sum_2397; // @[Mul.scala 207:34]
  wire  sum_2487 = cout_2394 ^ cout_2395; // @[Mul.scala 206:34]
  wire  cout_2487 = cout_2394 & cout_2395; // @[Mul.scala 207:34]
  wire  sum_2488 = sum_2398 ^ sum_2399; // @[Mul.scala 206:34]
  wire  cout_2488 = sum_2398 & sum_2399; // @[Mul.scala 207:34]
  wire  sum_2489 = cout_2396 ^ cout_2397; // @[Mul.scala 206:34]
  wire  cout_2489 = cout_2396 & cout_2397; // @[Mul.scala 207:34]
  wire  sum_2490 = sum_2400 ^ sum_2401; // @[Mul.scala 206:34]
  wire  cout_2490 = sum_2400 & sum_2401; // @[Mul.scala 207:34]
  wire  sum_2491 = cout_2398 ^ cout_2399; // @[Mul.scala 206:34]
  wire  cout_2491 = cout_2398 & cout_2399; // @[Mul.scala 207:34]
  wire  sum_2492 = sum_2402 ^ sum_2403; // @[Mul.scala 206:34]
  wire  cout_2492 = sum_2402 & sum_2403; // @[Mul.scala 207:34]
  wire  sum_2493 = cout_2400 ^ cout_2401; // @[Mul.scala 206:34]
  wire  cout_2493 = cout_2400 & cout_2401; // @[Mul.scala 207:34]
  wire  sum_2494 = sum_2404 ^ sum_2405; // @[Mul.scala 206:34]
  wire  cout_2494 = sum_2404 & sum_2405; // @[Mul.scala 207:34]
  wire  sum_2495 = cout_2402 ^ cout_2403; // @[Mul.scala 206:34]
  wire  cout_2495 = cout_2402 & cout_2403; // @[Mul.scala 207:34]
  wire  sum_2496 = sum_2406 ^ sum_2407; // @[Mul.scala 206:34]
  wire  cout_2496 = sum_2406 & sum_2407; // @[Mul.scala 207:34]
  wire  sum_2497 = cout_2404 ^ cout_2405; // @[Mul.scala 206:34]
  wire  cout_2497 = cout_2404 & cout_2405; // @[Mul.scala 207:34]
  wire  sum_2498 = sum_2408 ^ sum_2409; // @[Mul.scala 206:34]
  wire  cout_2498 = sum_2408 & sum_2409; // @[Mul.scala 207:34]
  wire  sum_2499 = cout_2406 ^ cout_2407; // @[Mul.scala 206:34]
  wire  cout_2499 = cout_2406 & cout_2407; // @[Mul.scala 207:34]
  wire  sum_2500 = sum_2410 ^ sum_2411; // @[Mul.scala 206:34]
  wire  cout_2500 = sum_2410 & sum_2411; // @[Mul.scala 207:34]
  wire  sum_2501 = cout_2408 ^ cout_2409; // @[Mul.scala 206:34]
  wire  cout_2501 = cout_2408 & cout_2409; // @[Mul.scala 207:34]
  wire  sum_2502 = sum_2412 ^ sum_2413; // @[Mul.scala 206:34]
  wire  cout_2502 = sum_2412 & sum_2413; // @[Mul.scala 207:34]
  wire  sum_2503 = cout_2410 ^ cout_2411; // @[Mul.scala 206:34]
  wire  cout_2503 = cout_2410 & cout_2411; // @[Mul.scala 207:34]
  wire  sum_2504 = sum_2414 ^ sum_2415; // @[Mul.scala 206:34]
  wire  cout_2504 = sum_2414 & sum_2415; // @[Mul.scala 207:34]
  wire  sum_2505 = cout_2412 ^ cout_2413; // @[Mul.scala 206:34]
  wire  cout_2505 = cout_2412 & cout_2413; // @[Mul.scala 207:34]
  wire  sum_2506 = sum_2416 ^ sum_2417; // @[Mul.scala 206:34]
  wire  cout_2506 = sum_2416 & sum_2417; // @[Mul.scala 207:34]
  wire  sum_2507 = cout_2414 ^ cout_2415; // @[Mul.scala 206:34]
  wire  cout_2507 = cout_2414 & cout_2415; // @[Mul.scala 207:34]
  wire  sum_2508 = sum_2418 ^ sum_2419; // @[Mul.scala 206:34]
  wire  cout_2508 = sum_2418 & sum_2419; // @[Mul.scala 207:34]
  wire  sum_2509 = cout_2416 ^ cout_2417; // @[Mul.scala 206:34]
  wire  cout_2509 = cout_2416 & cout_2417; // @[Mul.scala 207:34]
  wire  sum_2510 = sum_2420 ^ sum_2421; // @[Mul.scala 206:34]
  wire  cout_2510 = sum_2420 & sum_2421; // @[Mul.scala 207:34]
  wire  sum_2511 = cout_2418 ^ cout_2419; // @[Mul.scala 206:34]
  wire  cout_2511 = cout_2418 & cout_2419; // @[Mul.scala 207:34]
  wire  sum_2512 = sum_2422 ^ sum_2423; // @[Mul.scala 206:34]
  wire  cout_2512 = sum_2422 & sum_2423; // @[Mul.scala 207:34]
  wire  sum_2513 = cout_2420 ^ cout_2421; // @[Mul.scala 206:34]
  wire  cout_2513 = cout_2420 & cout_2421; // @[Mul.scala 207:34]
  wire  sum_2514 = sum_2424 ^ sum_2425; // @[Mul.scala 206:34]
  wire  cout_2514 = sum_2424 & sum_2425; // @[Mul.scala 207:34]
  wire  sum_2515 = cout_2422 ^ cout_2423; // @[Mul.scala 206:34]
  wire  cout_2515 = cout_2422 & cout_2423; // @[Mul.scala 207:34]
  wire  sum_2516 = sum_2426 ^ sum_2427; // @[Mul.scala 206:34]
  wire  cout_2516 = sum_2426 & sum_2427; // @[Mul.scala 207:34]
  wire  sum_2517 = cout_2424 ^ cout_2425; // @[Mul.scala 206:34]
  wire  cout_2517 = cout_2424 & cout_2425; // @[Mul.scala 207:34]
  wire  sum_2518 = sum_2428 ^ sum_2429; // @[Mul.scala 206:34]
  wire  cout_2518 = sum_2428 & sum_2429; // @[Mul.scala 207:34]
  wire  sum_2519 = cout_2426 ^ cout_2427; // @[Mul.scala 206:34]
  wire  cout_2519 = cout_2426 & cout_2427; // @[Mul.scala 207:34]
  wire  _sum_T_3170 = sum_2430 ^ cout_2428; // @[Mul.scala 191:34]
  wire  sum_2520 = sum_2430 ^ cout_2428 ^ cout_2429; // @[Mul.scala 191:42]
  wire  cout_2520 = sum_2430 & cout_2428 | _sum_T_3170 & cout_2429; // @[Mul.scala 192:44]
  wire  sum_2521 = sum_2431 ^ cout_2430; // @[Mul.scala 206:34]
  wire  cout_2521 = sum_2431 & cout_2430; // @[Mul.scala 207:34]
  wire  sum_2522 = sum_2432 ^ cout_2431; // @[Mul.scala 206:34]
  wire  cout_2522 = sum_2432 & cout_2431; // @[Mul.scala 207:34]
  wire  sum_2523 = sum_2433 ^ cout_2432; // @[Mul.scala 206:34]
  wire  cout_2523 = sum_2433 & cout_2432; // @[Mul.scala 207:34]
  wire  sum_2524 = sum_2434 ^ cout_2433; // @[Mul.scala 206:34]
  wire  cout_2524 = sum_2434 & cout_2433; // @[Mul.scala 207:34]
  wire  sum_2525 = sum_2435 ^ cout_2434; // @[Mul.scala 206:34]
  wire  sum_2553 = sum_2463 ^ cout_2462; // @[Mul.scala 206:34]
  wire  cout_2553 = sum_2463 & cout_2462; // @[Mul.scala 207:34]
  wire  sum_2554 = sum_2464 ^ cout_2463; // @[Mul.scala 206:34]
  wire  cout_2554 = sum_2464 & cout_2463; // @[Mul.scala 207:34]
  wire  sum_2555 = sum_2465 ^ cout_2464; // @[Mul.scala 206:34]
  wire  cout_2555 = sum_2465 & cout_2464; // @[Mul.scala 207:34]
  wire  _sum_T_3207 = sum_2466 ^ sum_2467; // @[Mul.scala 191:34]
  wire  sum_2556 = sum_2466 ^ sum_2467 ^ cout_2465; // @[Mul.scala 191:42]
  wire  cout_2556 = sum_2466 & sum_2467 | _sum_T_3207 & cout_2465; // @[Mul.scala 192:44]
  wire  sum_2557 = sum_2468 ^ sum_2469; // @[Mul.scala 206:34]
  wire  cout_2557 = sum_2468 & sum_2469; // @[Mul.scala 207:34]
  wire  sum_2558 = cout_2466 ^ cout_2467; // @[Mul.scala 206:34]
  wire  cout_2558 = cout_2466 & cout_2467; // @[Mul.scala 207:34]
  wire  sum_2559 = sum_2470 ^ sum_2471; // @[Mul.scala 206:34]
  wire  cout_2559 = sum_2470 & sum_2471; // @[Mul.scala 207:34]
  wire  sum_2560 = cout_2468 ^ cout_2469; // @[Mul.scala 206:34]
  wire  cout_2560 = cout_2468 & cout_2469; // @[Mul.scala 207:34]
  wire  sum_2561 = sum_2472 ^ sum_2473; // @[Mul.scala 206:34]
  wire  cout_2561 = sum_2472 & sum_2473; // @[Mul.scala 207:34]
  wire  sum_2562 = cout_2470 ^ cout_2471; // @[Mul.scala 206:34]
  wire  cout_2562 = cout_2470 & cout_2471; // @[Mul.scala 207:34]
  wire  sum_2563 = sum_2474 ^ sum_2475; // @[Mul.scala 206:34]
  wire  cout_2563 = sum_2474 & sum_2475; // @[Mul.scala 207:34]
  wire  sum_2564 = cout_2472 ^ cout_2473; // @[Mul.scala 206:34]
  wire  cout_2564 = cout_2472 & cout_2473; // @[Mul.scala 207:34]
  wire  sum_2565 = sum_2476 ^ sum_2477; // @[Mul.scala 206:34]
  wire  cout_2565 = sum_2476 & sum_2477; // @[Mul.scala 207:34]
  wire  sum_2566 = cout_2474 ^ cout_2475; // @[Mul.scala 206:34]
  wire  cout_2566 = cout_2474 & cout_2475; // @[Mul.scala 207:34]
  wire  sum_2567 = sum_2478 ^ sum_2479; // @[Mul.scala 206:34]
  wire  cout_2567 = sum_2478 & sum_2479; // @[Mul.scala 207:34]
  wire  sum_2568 = cout_2476 ^ cout_2477; // @[Mul.scala 206:34]
  wire  cout_2568 = cout_2476 & cout_2477; // @[Mul.scala 207:34]
  wire  sum_2569 = sum_2480 ^ sum_2481; // @[Mul.scala 206:34]
  wire  cout_2569 = sum_2480 & sum_2481; // @[Mul.scala 207:34]
  wire  sum_2570 = cout_2478 ^ cout_2479; // @[Mul.scala 206:34]
  wire  cout_2570 = cout_2478 & cout_2479; // @[Mul.scala 207:34]
  wire  sum_2571 = sum_2482 ^ sum_2483; // @[Mul.scala 206:34]
  wire  cout_2571 = sum_2482 & sum_2483; // @[Mul.scala 207:34]
  wire  sum_2572 = cout_2480 ^ cout_2481; // @[Mul.scala 206:34]
  wire  cout_2572 = cout_2480 & cout_2481; // @[Mul.scala 207:34]
  wire  sum_2573 = sum_2484 ^ sum_2485; // @[Mul.scala 206:34]
  wire  cout_2573 = sum_2484 & sum_2485; // @[Mul.scala 207:34]
  wire  sum_2574 = cout_2482 ^ cout_2483; // @[Mul.scala 206:34]
  wire  cout_2574 = cout_2482 & cout_2483; // @[Mul.scala 207:34]
  wire  sum_2575 = sum_2486 ^ sum_2487; // @[Mul.scala 206:34]
  wire  cout_2575 = sum_2486 & sum_2487; // @[Mul.scala 207:34]
  wire  sum_2576 = cout_2484 ^ cout_2485; // @[Mul.scala 206:34]
  wire  cout_2576 = cout_2484 & cout_2485; // @[Mul.scala 207:34]
  wire  sum_2577 = sum_2488 ^ sum_2489; // @[Mul.scala 206:34]
  wire  cout_2577 = sum_2488 & sum_2489; // @[Mul.scala 207:34]
  wire  sum_2578 = cout_2486 ^ cout_2487; // @[Mul.scala 206:34]
  wire  cout_2578 = cout_2486 & cout_2487; // @[Mul.scala 207:34]
  wire  sum_2579 = sum_2490 ^ sum_2491; // @[Mul.scala 206:34]
  wire  cout_2579 = sum_2490 & sum_2491; // @[Mul.scala 207:34]
  wire  sum_2580 = cout_2488 ^ cout_2489; // @[Mul.scala 206:34]
  wire  cout_2580 = cout_2488 & cout_2489; // @[Mul.scala 207:34]
  wire  sum_2581 = sum_2492 ^ sum_2493; // @[Mul.scala 206:34]
  wire  cout_2581 = sum_2492 & sum_2493; // @[Mul.scala 207:34]
  wire  sum_2582 = cout_2490 ^ cout_2491; // @[Mul.scala 206:34]
  wire  cout_2582 = cout_2490 & cout_2491; // @[Mul.scala 207:34]
  wire  sum_2583 = sum_2494 ^ sum_2495; // @[Mul.scala 206:34]
  wire  cout_2583 = sum_2494 & sum_2495; // @[Mul.scala 207:34]
  wire  sum_2584 = cout_2492 ^ cout_2493; // @[Mul.scala 206:34]
  wire  cout_2584 = cout_2492 & cout_2493; // @[Mul.scala 207:34]
  wire  sum_2585 = sum_2496 ^ sum_2497; // @[Mul.scala 206:34]
  wire  cout_2585 = sum_2496 & sum_2497; // @[Mul.scala 207:34]
  wire  sum_2586 = cout_2494 ^ cout_2495; // @[Mul.scala 206:34]
  wire  cout_2586 = cout_2494 & cout_2495; // @[Mul.scala 207:34]
  wire  sum_2587 = sum_2498 ^ sum_2499; // @[Mul.scala 206:34]
  wire  cout_2587 = sum_2498 & sum_2499; // @[Mul.scala 207:34]
  wire  sum_2588 = cout_2496 ^ cout_2497; // @[Mul.scala 206:34]
  wire  cout_2588 = cout_2496 & cout_2497; // @[Mul.scala 207:34]
  wire  sum_2589 = sum_2500 ^ sum_2501; // @[Mul.scala 206:34]
  wire  cout_2589 = sum_2500 & sum_2501; // @[Mul.scala 207:34]
  wire  sum_2590 = cout_2498 ^ cout_2499; // @[Mul.scala 206:34]
  wire  cout_2590 = cout_2498 & cout_2499; // @[Mul.scala 207:34]
  wire  sum_2591 = sum_2502 ^ sum_2503; // @[Mul.scala 206:34]
  wire  cout_2591 = sum_2502 & sum_2503; // @[Mul.scala 207:34]
  wire  sum_2592 = cout_2500 ^ cout_2501; // @[Mul.scala 206:34]
  wire  cout_2592 = cout_2500 & cout_2501; // @[Mul.scala 207:34]
  wire  sum_2593 = sum_2504 ^ sum_2505; // @[Mul.scala 206:34]
  wire  cout_2593 = sum_2504 & sum_2505; // @[Mul.scala 207:34]
  wire  sum_2594 = cout_2502 ^ cout_2503; // @[Mul.scala 206:34]
  wire  cout_2594 = cout_2502 & cout_2503; // @[Mul.scala 207:34]
  wire  sum_2595 = sum_2506 ^ sum_2507; // @[Mul.scala 206:34]
  wire  cout_2595 = sum_2506 & sum_2507; // @[Mul.scala 207:34]
  wire  sum_2596 = cout_2504 ^ cout_2505; // @[Mul.scala 206:34]
  wire  cout_2596 = cout_2504 & cout_2505; // @[Mul.scala 207:34]
  wire  sum_2597 = sum_2508 ^ sum_2509; // @[Mul.scala 206:34]
  wire  cout_2597 = sum_2508 & sum_2509; // @[Mul.scala 207:34]
  wire  sum_2598 = cout_2506 ^ cout_2507; // @[Mul.scala 206:34]
  wire  cout_2598 = cout_2506 & cout_2507; // @[Mul.scala 207:34]
  wire  sum_2599 = sum_2510 ^ sum_2511; // @[Mul.scala 206:34]
  wire  cout_2599 = sum_2510 & sum_2511; // @[Mul.scala 207:34]
  wire  sum_2600 = cout_2508 ^ cout_2509; // @[Mul.scala 206:34]
  wire  cout_2600 = cout_2508 & cout_2509; // @[Mul.scala 207:34]
  wire  sum_2601 = sum_2512 ^ sum_2513; // @[Mul.scala 206:34]
  wire  cout_2601 = sum_2512 & sum_2513; // @[Mul.scala 207:34]
  wire  sum_2602 = cout_2510 ^ cout_2511; // @[Mul.scala 206:34]
  wire  cout_2602 = cout_2510 & cout_2511; // @[Mul.scala 207:34]
  wire  sum_2603 = sum_2514 ^ sum_2515; // @[Mul.scala 206:34]
  wire  cout_2603 = sum_2514 & sum_2515; // @[Mul.scala 207:34]
  wire  sum_2604 = cout_2512 ^ cout_2513; // @[Mul.scala 206:34]
  wire  cout_2604 = cout_2512 & cout_2513; // @[Mul.scala 207:34]
  wire  sum_2605 = sum_2516 ^ sum_2517; // @[Mul.scala 206:34]
  wire  cout_2605 = sum_2516 & sum_2517; // @[Mul.scala 207:34]
  wire  sum_2606 = cout_2514 ^ cout_2515; // @[Mul.scala 206:34]
  wire  cout_2606 = cout_2514 & cout_2515; // @[Mul.scala 207:34]
  wire  sum_2607 = sum_2518 ^ sum_2519; // @[Mul.scala 206:34]
  wire  cout_2607 = sum_2518 & sum_2519; // @[Mul.scala 207:34]
  wire  sum_2608 = cout_2516 ^ cout_2517; // @[Mul.scala 206:34]
  wire  cout_2608 = cout_2516 & cout_2517; // @[Mul.scala 207:34]
  wire  _sum_T_3261 = sum_2520 ^ cout_2518; // @[Mul.scala 191:34]
  wire  sum_2609 = sum_2520 ^ cout_2518 ^ cout_2519; // @[Mul.scala 191:42]
  wire  cout_2609 = sum_2520 & cout_2518 | _sum_T_3261 & cout_2519; // @[Mul.scala 192:44]
  wire  sum_2610 = sum_2521 ^ cout_2520; // @[Mul.scala 206:34]
  wire  cout_2610 = sum_2521 & cout_2520; // @[Mul.scala 207:34]
  wire  sum_2611 = sum_2522 ^ cout_2521; // @[Mul.scala 206:34]
  wire  cout_2611 = sum_2522 & cout_2521; // @[Mul.scala 207:34]
  wire  sum_2612 = sum_2523 ^ cout_2522; // @[Mul.scala 206:34]
  wire  cout_2612 = sum_2523 & cout_2522; // @[Mul.scala 207:34]
  wire  sum_2613 = sum_2524 ^ cout_2523; // @[Mul.scala 206:34]
  wire  cout_2613 = sum_2524 & cout_2523; // @[Mul.scala 207:34]
  wire  sum_2614 = sum_2525 ^ cout_2524; // @[Mul.scala 206:34]
  wire  sum_2643 = sum_2554 ^ cout_2553; // @[Mul.scala 206:34]
  wire  cout_2643 = sum_2554 & cout_2553; // @[Mul.scala 207:34]
  wire  sum_2644 = sum_2555 ^ cout_2554; // @[Mul.scala 206:34]
  wire  cout_2644 = sum_2555 & cout_2554; // @[Mul.scala 207:34]
  wire  sum_2645 = sum_2556 ^ cout_2555; // @[Mul.scala 206:34]
  wire  cout_2645 = sum_2556 & cout_2555; // @[Mul.scala 207:34]
  wire  _sum_T_3299 = sum_2557 ^ sum_2558; // @[Mul.scala 191:34]
  wire  sum_2646 = sum_2557 ^ sum_2558 ^ cout_2556; // @[Mul.scala 191:42]
  wire  cout_2646 = sum_2557 & sum_2558 | _sum_T_3299 & cout_2556; // @[Mul.scala 192:44]
  wire  sum_2647 = sum_2559 ^ sum_2560; // @[Mul.scala 206:34]
  wire  cout_2647 = sum_2559 & sum_2560; // @[Mul.scala 207:34]
  wire  sum_2648 = cout_2557 ^ cout_2558; // @[Mul.scala 206:34]
  wire  cout_2648 = cout_2557 & cout_2558; // @[Mul.scala 207:34]
  wire  sum_2649 = sum_2561 ^ sum_2562; // @[Mul.scala 206:34]
  wire  cout_2649 = sum_2561 & sum_2562; // @[Mul.scala 207:34]
  wire  sum_2650 = cout_2559 ^ cout_2560; // @[Mul.scala 206:34]
  wire  cout_2650 = cout_2559 & cout_2560; // @[Mul.scala 207:34]
  wire  sum_2651 = sum_2563 ^ sum_2564; // @[Mul.scala 206:34]
  wire  cout_2651 = sum_2563 & sum_2564; // @[Mul.scala 207:34]
  wire  sum_2652 = cout_2561 ^ cout_2562; // @[Mul.scala 206:34]
  wire  cout_2652 = cout_2561 & cout_2562; // @[Mul.scala 207:34]
  wire  sum_2653 = sum_2565 ^ sum_2566; // @[Mul.scala 206:34]
  wire  cout_2653 = sum_2565 & sum_2566; // @[Mul.scala 207:34]
  wire  sum_2654 = cout_2563 ^ cout_2564; // @[Mul.scala 206:34]
  wire  cout_2654 = cout_2563 & cout_2564; // @[Mul.scala 207:34]
  wire  sum_2655 = sum_2567 ^ sum_2568; // @[Mul.scala 206:34]
  wire  cout_2655 = sum_2567 & sum_2568; // @[Mul.scala 207:34]
  wire  sum_2656 = cout_2565 ^ cout_2566; // @[Mul.scala 206:34]
  wire  cout_2656 = cout_2565 & cout_2566; // @[Mul.scala 207:34]
  wire  sum_2657 = sum_2569 ^ sum_2570; // @[Mul.scala 206:34]
  wire  cout_2657 = sum_2569 & sum_2570; // @[Mul.scala 207:34]
  wire  sum_2658 = cout_2567 ^ cout_2568; // @[Mul.scala 206:34]
  wire  cout_2658 = cout_2567 & cout_2568; // @[Mul.scala 207:34]
  wire  sum_2659 = sum_2571 ^ sum_2572; // @[Mul.scala 206:34]
  wire  cout_2659 = sum_2571 & sum_2572; // @[Mul.scala 207:34]
  wire  sum_2660 = cout_2569 ^ cout_2570; // @[Mul.scala 206:34]
  wire  cout_2660 = cout_2569 & cout_2570; // @[Mul.scala 207:34]
  wire  sum_2661 = sum_2573 ^ sum_2574; // @[Mul.scala 206:34]
  wire  cout_2661 = sum_2573 & sum_2574; // @[Mul.scala 207:34]
  wire  sum_2662 = cout_2571 ^ cout_2572; // @[Mul.scala 206:34]
  wire  cout_2662 = cout_2571 & cout_2572; // @[Mul.scala 207:34]
  wire  sum_2663 = sum_2575 ^ sum_2576; // @[Mul.scala 206:34]
  wire  cout_2663 = sum_2575 & sum_2576; // @[Mul.scala 207:34]
  wire  sum_2664 = cout_2573 ^ cout_2574; // @[Mul.scala 206:34]
  wire  cout_2664 = cout_2573 & cout_2574; // @[Mul.scala 207:34]
  wire  sum_2665 = sum_2577 ^ sum_2578; // @[Mul.scala 206:34]
  wire  cout_2665 = sum_2577 & sum_2578; // @[Mul.scala 207:34]
  wire  sum_2666 = cout_2575 ^ cout_2576; // @[Mul.scala 206:34]
  wire  cout_2666 = cout_2575 & cout_2576; // @[Mul.scala 207:34]
  wire  sum_2667 = sum_2579 ^ sum_2580; // @[Mul.scala 206:34]
  wire  cout_2667 = sum_2579 & sum_2580; // @[Mul.scala 207:34]
  wire  sum_2668 = cout_2577 ^ cout_2578; // @[Mul.scala 206:34]
  wire  cout_2668 = cout_2577 & cout_2578; // @[Mul.scala 207:34]
  wire  sum_2669 = sum_2581 ^ sum_2582; // @[Mul.scala 206:34]
  wire  cout_2669 = sum_2581 & sum_2582; // @[Mul.scala 207:34]
  wire  sum_2670 = cout_2579 ^ cout_2580; // @[Mul.scala 206:34]
  wire  cout_2670 = cout_2579 & cout_2580; // @[Mul.scala 207:34]
  wire  sum_2671 = sum_2583 ^ sum_2584; // @[Mul.scala 206:34]
  wire  cout_2671 = sum_2583 & sum_2584; // @[Mul.scala 207:34]
  wire  sum_2672 = cout_2581 ^ cout_2582; // @[Mul.scala 206:34]
  wire  cout_2672 = cout_2581 & cout_2582; // @[Mul.scala 207:34]
  wire  sum_2673 = sum_2585 ^ sum_2586; // @[Mul.scala 206:34]
  wire  cout_2673 = sum_2585 & sum_2586; // @[Mul.scala 207:34]
  wire  sum_2674 = cout_2583 ^ cout_2584; // @[Mul.scala 206:34]
  wire  cout_2674 = cout_2583 & cout_2584; // @[Mul.scala 207:34]
  wire  sum_2675 = sum_2587 ^ sum_2588; // @[Mul.scala 206:34]
  wire  cout_2675 = sum_2587 & sum_2588; // @[Mul.scala 207:34]
  wire  sum_2676 = cout_2585 ^ cout_2586; // @[Mul.scala 206:34]
  wire  cout_2676 = cout_2585 & cout_2586; // @[Mul.scala 207:34]
  wire  sum_2677 = sum_2589 ^ sum_2590; // @[Mul.scala 206:34]
  wire  cout_2677 = sum_2589 & sum_2590; // @[Mul.scala 207:34]
  wire  sum_2678 = cout_2587 ^ cout_2588; // @[Mul.scala 206:34]
  wire  cout_2678 = cout_2587 & cout_2588; // @[Mul.scala 207:34]
  wire  sum_2679 = sum_2591 ^ sum_2592; // @[Mul.scala 206:34]
  wire  cout_2679 = sum_2591 & sum_2592; // @[Mul.scala 207:34]
  wire  sum_2680 = cout_2589 ^ cout_2590; // @[Mul.scala 206:34]
  wire  cout_2680 = cout_2589 & cout_2590; // @[Mul.scala 207:34]
  wire  sum_2681 = sum_2593 ^ sum_2594; // @[Mul.scala 206:34]
  wire  cout_2681 = sum_2593 & sum_2594; // @[Mul.scala 207:34]
  wire  sum_2682 = cout_2591 ^ cout_2592; // @[Mul.scala 206:34]
  wire  cout_2682 = cout_2591 & cout_2592; // @[Mul.scala 207:34]
  wire  sum_2683 = sum_2595 ^ sum_2596; // @[Mul.scala 206:34]
  wire  cout_2683 = sum_2595 & sum_2596; // @[Mul.scala 207:34]
  wire  sum_2684 = cout_2593 ^ cout_2594; // @[Mul.scala 206:34]
  wire  cout_2684 = cout_2593 & cout_2594; // @[Mul.scala 207:34]
  wire  sum_2685 = sum_2597 ^ sum_2598; // @[Mul.scala 206:34]
  wire  cout_2685 = sum_2597 & sum_2598; // @[Mul.scala 207:34]
  wire  sum_2686 = cout_2595 ^ cout_2596; // @[Mul.scala 206:34]
  wire  cout_2686 = cout_2595 & cout_2596; // @[Mul.scala 207:34]
  wire  sum_2687 = sum_2599 ^ sum_2600; // @[Mul.scala 206:34]
  wire  cout_2687 = sum_2599 & sum_2600; // @[Mul.scala 207:34]
  wire  sum_2688 = cout_2597 ^ cout_2598; // @[Mul.scala 206:34]
  wire  cout_2688 = cout_2597 & cout_2598; // @[Mul.scala 207:34]
  wire  sum_2689 = sum_2601 ^ sum_2602; // @[Mul.scala 206:34]
  wire  cout_2689 = sum_2601 & sum_2602; // @[Mul.scala 207:34]
  wire  sum_2690 = cout_2599 ^ cout_2600; // @[Mul.scala 206:34]
  wire  cout_2690 = cout_2599 & cout_2600; // @[Mul.scala 207:34]
  wire  sum_2691 = sum_2603 ^ sum_2604; // @[Mul.scala 206:34]
  wire  cout_2691 = sum_2603 & sum_2604; // @[Mul.scala 207:34]
  wire  sum_2692 = cout_2601 ^ cout_2602; // @[Mul.scala 206:34]
  wire  cout_2692 = cout_2601 & cout_2602; // @[Mul.scala 207:34]
  wire  sum_2693 = sum_2605 ^ sum_2606; // @[Mul.scala 206:34]
  wire  cout_2693 = sum_2605 & sum_2606; // @[Mul.scala 207:34]
  wire  sum_2694 = cout_2603 ^ cout_2604; // @[Mul.scala 206:34]
  wire  cout_2694 = cout_2603 & cout_2604; // @[Mul.scala 207:34]
  wire  sum_2695 = sum_2607 ^ sum_2608; // @[Mul.scala 206:34]
  wire  cout_2695 = sum_2607 & sum_2608; // @[Mul.scala 207:34]
  wire  sum_2696 = cout_2605 ^ cout_2606; // @[Mul.scala 206:34]
  wire  cout_2696 = cout_2605 & cout_2606; // @[Mul.scala 207:34]
  wire  _sum_T_3351 = sum_2609 ^ cout_2607; // @[Mul.scala 191:34]
  wire  sum_2697 = sum_2609 ^ cout_2607 ^ cout_2608; // @[Mul.scala 191:42]
  wire  cout_2697 = sum_2609 & cout_2607 | _sum_T_3351 & cout_2608; // @[Mul.scala 192:44]
  wire  sum_2698 = sum_2610 ^ cout_2609; // @[Mul.scala 206:34]
  wire  cout_2698 = sum_2610 & cout_2609; // @[Mul.scala 207:34]
  wire  sum_2699 = sum_2611 ^ cout_2610; // @[Mul.scala 206:34]
  wire  cout_2699 = sum_2611 & cout_2610; // @[Mul.scala 207:34]
  wire  sum_2700 = sum_2612 ^ cout_2611; // @[Mul.scala 206:34]
  wire  cout_2700 = sum_2612 & cout_2611; // @[Mul.scala 207:34]
  wire  sum_2701 = sum_2613 ^ cout_2612; // @[Mul.scala 206:34]
  wire  cout_2701 = sum_2613 & cout_2612; // @[Mul.scala 207:34]
  wire  sum_2702 = sum_2614 ^ cout_2613; // @[Mul.scala 206:34]
  wire  sum_2732 = sum_2644 ^ cout_2643; // @[Mul.scala 206:34]
  wire  cout_2732 = sum_2644 & cout_2643; // @[Mul.scala 207:34]
  wire  sum_2733 = sum_2645 ^ cout_2644; // @[Mul.scala 206:34]
  wire  cout_2733 = sum_2645 & cout_2644; // @[Mul.scala 207:34]
  wire  sum_2734 = sum_2646 ^ cout_2645; // @[Mul.scala 206:34]
  wire  cout_2734 = sum_2646 & cout_2645; // @[Mul.scala 207:34]
  wire  _sum_T_3390 = sum_2647 ^ sum_2648; // @[Mul.scala 191:34]
  wire  sum_2735 = sum_2647 ^ sum_2648 ^ cout_2646; // @[Mul.scala 191:42]
  wire  cout_2735 = sum_2647 & sum_2648 | _sum_T_3390 & cout_2646; // @[Mul.scala 192:44]
  wire  sum_2736 = sum_2649 ^ sum_2650; // @[Mul.scala 206:34]
  wire  cout_2736 = sum_2649 & sum_2650; // @[Mul.scala 207:34]
  wire  sum_2737 = cout_2647 ^ cout_2648; // @[Mul.scala 206:34]
  wire  cout_2737 = cout_2647 & cout_2648; // @[Mul.scala 207:34]
  wire  sum_2738 = sum_2651 ^ sum_2652; // @[Mul.scala 206:34]
  wire  cout_2738 = sum_2651 & sum_2652; // @[Mul.scala 207:34]
  wire  sum_2739 = cout_2649 ^ cout_2650; // @[Mul.scala 206:34]
  wire  cout_2739 = cout_2649 & cout_2650; // @[Mul.scala 207:34]
  wire  sum_2740 = sum_2653 ^ sum_2654; // @[Mul.scala 206:34]
  wire  cout_2740 = sum_2653 & sum_2654; // @[Mul.scala 207:34]
  wire  sum_2741 = cout_2651 ^ cout_2652; // @[Mul.scala 206:34]
  wire  cout_2741 = cout_2651 & cout_2652; // @[Mul.scala 207:34]
  wire  sum_2742 = sum_2655 ^ sum_2656; // @[Mul.scala 206:34]
  wire  cout_2742 = sum_2655 & sum_2656; // @[Mul.scala 207:34]
  wire  sum_2743 = cout_2653 ^ cout_2654; // @[Mul.scala 206:34]
  wire  cout_2743 = cout_2653 & cout_2654; // @[Mul.scala 207:34]
  wire  sum_2744 = sum_2657 ^ sum_2658; // @[Mul.scala 206:34]
  wire  cout_2744 = sum_2657 & sum_2658; // @[Mul.scala 207:34]
  wire  sum_2745 = cout_2655 ^ cout_2656; // @[Mul.scala 206:34]
  wire  cout_2745 = cout_2655 & cout_2656; // @[Mul.scala 207:34]
  wire  sum_2746 = sum_2659 ^ sum_2660; // @[Mul.scala 206:34]
  wire  cout_2746 = sum_2659 & sum_2660; // @[Mul.scala 207:34]
  wire  sum_2747 = cout_2657 ^ cout_2658; // @[Mul.scala 206:34]
  wire  cout_2747 = cout_2657 & cout_2658; // @[Mul.scala 207:34]
  wire  sum_2748 = sum_2661 ^ sum_2662; // @[Mul.scala 206:34]
  wire  cout_2748 = sum_2661 & sum_2662; // @[Mul.scala 207:34]
  wire  sum_2749 = cout_2659 ^ cout_2660; // @[Mul.scala 206:34]
  wire  cout_2749 = cout_2659 & cout_2660; // @[Mul.scala 207:34]
  wire  sum_2750 = sum_2663 ^ sum_2664; // @[Mul.scala 206:34]
  wire  cout_2750 = sum_2663 & sum_2664; // @[Mul.scala 207:34]
  wire  sum_2751 = cout_2661 ^ cout_2662; // @[Mul.scala 206:34]
  wire  cout_2751 = cout_2661 & cout_2662; // @[Mul.scala 207:34]
  wire  sum_2752 = sum_2665 ^ sum_2666; // @[Mul.scala 206:34]
  wire  cout_2752 = sum_2665 & sum_2666; // @[Mul.scala 207:34]
  wire  sum_2753 = cout_2663 ^ cout_2664; // @[Mul.scala 206:34]
  wire  cout_2753 = cout_2663 & cout_2664; // @[Mul.scala 207:34]
  wire  sum_2754 = sum_2667 ^ sum_2668; // @[Mul.scala 206:34]
  wire  cout_2754 = sum_2667 & sum_2668; // @[Mul.scala 207:34]
  wire  sum_2755 = cout_2665 ^ cout_2666; // @[Mul.scala 206:34]
  wire  cout_2755 = cout_2665 & cout_2666; // @[Mul.scala 207:34]
  wire  sum_2756 = sum_2669 ^ sum_2670; // @[Mul.scala 206:34]
  wire  cout_2756 = sum_2669 & sum_2670; // @[Mul.scala 207:34]
  wire  sum_2757 = cout_2667 ^ cout_2668; // @[Mul.scala 206:34]
  wire  cout_2757 = cout_2667 & cout_2668; // @[Mul.scala 207:34]
  wire  sum_2758 = sum_2671 ^ sum_2672; // @[Mul.scala 206:34]
  wire  cout_2758 = sum_2671 & sum_2672; // @[Mul.scala 207:34]
  wire  sum_2759 = cout_2669 ^ cout_2670; // @[Mul.scala 206:34]
  wire  cout_2759 = cout_2669 & cout_2670; // @[Mul.scala 207:34]
  wire  sum_2760 = sum_2673 ^ sum_2674; // @[Mul.scala 206:34]
  wire  cout_2760 = sum_2673 & sum_2674; // @[Mul.scala 207:34]
  wire  sum_2761 = cout_2671 ^ cout_2672; // @[Mul.scala 206:34]
  wire  cout_2761 = cout_2671 & cout_2672; // @[Mul.scala 207:34]
  wire  sum_2762 = sum_2675 ^ sum_2676; // @[Mul.scala 206:34]
  wire  cout_2762 = sum_2675 & sum_2676; // @[Mul.scala 207:34]
  wire  sum_2763 = cout_2673 ^ cout_2674; // @[Mul.scala 206:34]
  wire  cout_2763 = cout_2673 & cout_2674; // @[Mul.scala 207:34]
  wire  sum_2764 = sum_2677 ^ sum_2678; // @[Mul.scala 206:34]
  wire  cout_2764 = sum_2677 & sum_2678; // @[Mul.scala 207:34]
  wire  sum_2765 = cout_2675 ^ cout_2676; // @[Mul.scala 206:34]
  wire  cout_2765 = cout_2675 & cout_2676; // @[Mul.scala 207:34]
  wire  sum_2766 = sum_2679 ^ sum_2680; // @[Mul.scala 206:34]
  wire  cout_2766 = sum_2679 & sum_2680; // @[Mul.scala 207:34]
  wire  sum_2767 = cout_2677 ^ cout_2678; // @[Mul.scala 206:34]
  wire  cout_2767 = cout_2677 & cout_2678; // @[Mul.scala 207:34]
  wire  sum_2768 = sum_2681 ^ sum_2682; // @[Mul.scala 206:34]
  wire  cout_2768 = sum_2681 & sum_2682; // @[Mul.scala 207:34]
  wire  sum_2769 = cout_2679 ^ cout_2680; // @[Mul.scala 206:34]
  wire  cout_2769 = cout_2679 & cout_2680; // @[Mul.scala 207:34]
  wire  sum_2770 = sum_2683 ^ sum_2684; // @[Mul.scala 206:34]
  wire  cout_2770 = sum_2683 & sum_2684; // @[Mul.scala 207:34]
  wire  sum_2771 = cout_2681 ^ cout_2682; // @[Mul.scala 206:34]
  wire  cout_2771 = cout_2681 & cout_2682; // @[Mul.scala 207:34]
  wire  sum_2772 = sum_2685 ^ sum_2686; // @[Mul.scala 206:34]
  wire  cout_2772 = sum_2685 & sum_2686; // @[Mul.scala 207:34]
  wire  sum_2773 = cout_2683 ^ cout_2684; // @[Mul.scala 206:34]
  wire  cout_2773 = cout_2683 & cout_2684; // @[Mul.scala 207:34]
  wire  sum_2774 = sum_2687 ^ sum_2688; // @[Mul.scala 206:34]
  wire  cout_2774 = sum_2687 & sum_2688; // @[Mul.scala 207:34]
  wire  sum_2775 = cout_2685 ^ cout_2686; // @[Mul.scala 206:34]
  wire  cout_2775 = cout_2685 & cout_2686; // @[Mul.scala 207:34]
  wire  sum_2776 = sum_2689 ^ sum_2690; // @[Mul.scala 206:34]
  wire  cout_2776 = sum_2689 & sum_2690; // @[Mul.scala 207:34]
  wire  sum_2777 = cout_2687 ^ cout_2688; // @[Mul.scala 206:34]
  wire  cout_2777 = cout_2687 & cout_2688; // @[Mul.scala 207:34]
  wire  sum_2778 = sum_2691 ^ sum_2692; // @[Mul.scala 206:34]
  wire  cout_2778 = sum_2691 & sum_2692; // @[Mul.scala 207:34]
  wire  sum_2779 = cout_2689 ^ cout_2690; // @[Mul.scala 206:34]
  wire  cout_2779 = cout_2689 & cout_2690; // @[Mul.scala 207:34]
  wire  sum_2780 = sum_2693 ^ sum_2694; // @[Mul.scala 206:34]
  wire  cout_2780 = sum_2693 & sum_2694; // @[Mul.scala 207:34]
  wire  sum_2781 = cout_2691 ^ cout_2692; // @[Mul.scala 206:34]
  wire  cout_2781 = cout_2691 & cout_2692; // @[Mul.scala 207:34]
  wire  sum_2782 = sum_2695 ^ sum_2696; // @[Mul.scala 206:34]
  wire  cout_2782 = sum_2695 & sum_2696; // @[Mul.scala 207:34]
  wire  sum_2783 = cout_2693 ^ cout_2694; // @[Mul.scala 206:34]
  wire  cout_2783 = cout_2693 & cout_2694; // @[Mul.scala 207:34]
  wire  _sum_T_3440 = sum_2697 ^ cout_2695; // @[Mul.scala 191:34]
  wire  sum_2784 = sum_2697 ^ cout_2695 ^ cout_2696; // @[Mul.scala 191:42]
  wire  cout_2784 = sum_2697 & cout_2695 | _sum_T_3440 & cout_2696; // @[Mul.scala 192:44]
  wire  sum_2785 = sum_2698 ^ cout_2697; // @[Mul.scala 206:34]
  wire  cout_2785 = sum_2698 & cout_2697; // @[Mul.scala 207:34]
  wire  sum_2786 = sum_2699 ^ cout_2698; // @[Mul.scala 206:34]
  wire  cout_2786 = sum_2699 & cout_2698; // @[Mul.scala 207:34]
  wire  sum_2787 = sum_2700 ^ cout_2699; // @[Mul.scala 206:34]
  wire  cout_2787 = sum_2700 & cout_2699; // @[Mul.scala 207:34]
  wire  sum_2788 = sum_2701 ^ cout_2700; // @[Mul.scala 206:34]
  wire  cout_2788 = sum_2701 & cout_2700; // @[Mul.scala 207:34]
  wire  sum_2789 = sum_2702 ^ cout_2701; // @[Mul.scala 206:34]
  wire  sum_2820 = sum_2733 ^ cout_2732; // @[Mul.scala 206:34]
  wire  cout_2820 = sum_2733 & cout_2732; // @[Mul.scala 207:34]
  wire  sum_2821 = sum_2734 ^ cout_2733; // @[Mul.scala 206:34]
  wire  cout_2821 = sum_2734 & cout_2733; // @[Mul.scala 207:34]
  wire  sum_2822 = sum_2735 ^ cout_2734; // @[Mul.scala 206:34]
  wire  cout_2822 = sum_2735 & cout_2734; // @[Mul.scala 207:34]
  wire  _sum_T_3480 = sum_2736 ^ sum_2737; // @[Mul.scala 191:34]
  wire  sum_2823 = sum_2736 ^ sum_2737 ^ cout_2735; // @[Mul.scala 191:42]
  wire  cout_2823 = sum_2736 & sum_2737 | _sum_T_3480 & cout_2735; // @[Mul.scala 192:44]
  wire  sum_2824 = sum_2738 ^ sum_2739; // @[Mul.scala 206:34]
  wire  cout_2824 = sum_2738 & sum_2739; // @[Mul.scala 207:34]
  wire  sum_2825 = cout_2736 ^ cout_2737; // @[Mul.scala 206:34]
  wire  cout_2825 = cout_2736 & cout_2737; // @[Mul.scala 207:34]
  wire  sum_2826 = sum_2740 ^ sum_2741; // @[Mul.scala 206:34]
  wire  cout_2826 = sum_2740 & sum_2741; // @[Mul.scala 207:34]
  wire  sum_2827 = cout_2738 ^ cout_2739; // @[Mul.scala 206:34]
  wire  cout_2827 = cout_2738 & cout_2739; // @[Mul.scala 207:34]
  wire  sum_2828 = sum_2742 ^ sum_2743; // @[Mul.scala 206:34]
  wire  cout_2828 = sum_2742 & sum_2743; // @[Mul.scala 207:34]
  wire  sum_2829 = cout_2740 ^ cout_2741; // @[Mul.scala 206:34]
  wire  cout_2829 = cout_2740 & cout_2741; // @[Mul.scala 207:34]
  wire  sum_2830 = sum_2744 ^ sum_2745; // @[Mul.scala 206:34]
  wire  cout_2830 = sum_2744 & sum_2745; // @[Mul.scala 207:34]
  wire  sum_2831 = cout_2742 ^ cout_2743; // @[Mul.scala 206:34]
  wire  cout_2831 = cout_2742 & cout_2743; // @[Mul.scala 207:34]
  wire  sum_2832 = sum_2746 ^ sum_2747; // @[Mul.scala 206:34]
  wire  cout_2832 = sum_2746 & sum_2747; // @[Mul.scala 207:34]
  wire  sum_2833 = cout_2744 ^ cout_2745; // @[Mul.scala 206:34]
  wire  cout_2833 = cout_2744 & cout_2745; // @[Mul.scala 207:34]
  wire  sum_2834 = sum_2748 ^ sum_2749; // @[Mul.scala 206:34]
  wire  cout_2834 = sum_2748 & sum_2749; // @[Mul.scala 207:34]
  wire  sum_2835 = cout_2746 ^ cout_2747; // @[Mul.scala 206:34]
  wire  cout_2835 = cout_2746 & cout_2747; // @[Mul.scala 207:34]
  wire  sum_2836 = sum_2750 ^ sum_2751; // @[Mul.scala 206:34]
  wire  cout_2836 = sum_2750 & sum_2751; // @[Mul.scala 207:34]
  wire  sum_2837 = cout_2748 ^ cout_2749; // @[Mul.scala 206:34]
  wire  cout_2837 = cout_2748 & cout_2749; // @[Mul.scala 207:34]
  wire  sum_2838 = sum_2752 ^ sum_2753; // @[Mul.scala 206:34]
  wire  cout_2838 = sum_2752 & sum_2753; // @[Mul.scala 207:34]
  wire  sum_2839 = cout_2750 ^ cout_2751; // @[Mul.scala 206:34]
  wire  cout_2839 = cout_2750 & cout_2751; // @[Mul.scala 207:34]
  wire  sum_2840 = sum_2754 ^ sum_2755; // @[Mul.scala 206:34]
  wire  cout_2840 = sum_2754 & sum_2755; // @[Mul.scala 207:34]
  wire  sum_2841 = cout_2752 ^ cout_2753; // @[Mul.scala 206:34]
  wire  cout_2841 = cout_2752 & cout_2753; // @[Mul.scala 207:34]
  wire  sum_2842 = sum_2756 ^ sum_2757; // @[Mul.scala 206:34]
  wire  cout_2842 = sum_2756 & sum_2757; // @[Mul.scala 207:34]
  wire  sum_2843 = cout_2754 ^ cout_2755; // @[Mul.scala 206:34]
  wire  cout_2843 = cout_2754 & cout_2755; // @[Mul.scala 207:34]
  wire  sum_2844 = sum_2758 ^ sum_2759; // @[Mul.scala 206:34]
  wire  cout_2844 = sum_2758 & sum_2759; // @[Mul.scala 207:34]
  wire  sum_2845 = cout_2756 ^ cout_2757; // @[Mul.scala 206:34]
  wire  cout_2845 = cout_2756 & cout_2757; // @[Mul.scala 207:34]
  wire  sum_2846 = sum_2760 ^ sum_2761; // @[Mul.scala 206:34]
  wire  cout_2846 = sum_2760 & sum_2761; // @[Mul.scala 207:34]
  wire  sum_2847 = cout_2758 ^ cout_2759; // @[Mul.scala 206:34]
  wire  cout_2847 = cout_2758 & cout_2759; // @[Mul.scala 207:34]
  wire  sum_2848 = sum_2762 ^ sum_2763; // @[Mul.scala 206:34]
  wire  cout_2848 = sum_2762 & sum_2763; // @[Mul.scala 207:34]
  wire  sum_2849 = cout_2760 ^ cout_2761; // @[Mul.scala 206:34]
  wire  cout_2849 = cout_2760 & cout_2761; // @[Mul.scala 207:34]
  wire  sum_2850 = sum_2764 ^ sum_2765; // @[Mul.scala 206:34]
  wire  cout_2850 = sum_2764 & sum_2765; // @[Mul.scala 207:34]
  wire  sum_2851 = cout_2762 ^ cout_2763; // @[Mul.scala 206:34]
  wire  cout_2851 = cout_2762 & cout_2763; // @[Mul.scala 207:34]
  wire  sum_2852 = sum_2766 ^ sum_2767; // @[Mul.scala 206:34]
  wire  cout_2852 = sum_2766 & sum_2767; // @[Mul.scala 207:34]
  wire  sum_2853 = cout_2764 ^ cout_2765; // @[Mul.scala 206:34]
  wire  cout_2853 = cout_2764 & cout_2765; // @[Mul.scala 207:34]
  wire  sum_2854 = sum_2768 ^ sum_2769; // @[Mul.scala 206:34]
  wire  cout_2854 = sum_2768 & sum_2769; // @[Mul.scala 207:34]
  wire  sum_2855 = cout_2766 ^ cout_2767; // @[Mul.scala 206:34]
  wire  cout_2855 = cout_2766 & cout_2767; // @[Mul.scala 207:34]
  wire  sum_2856 = sum_2770 ^ sum_2771; // @[Mul.scala 206:34]
  wire  cout_2856 = sum_2770 & sum_2771; // @[Mul.scala 207:34]
  wire  sum_2857 = cout_2768 ^ cout_2769; // @[Mul.scala 206:34]
  wire  cout_2857 = cout_2768 & cout_2769; // @[Mul.scala 207:34]
  wire  sum_2858 = sum_2772 ^ sum_2773; // @[Mul.scala 206:34]
  wire  cout_2858 = sum_2772 & sum_2773; // @[Mul.scala 207:34]
  wire  sum_2859 = cout_2770 ^ cout_2771; // @[Mul.scala 206:34]
  wire  cout_2859 = cout_2770 & cout_2771; // @[Mul.scala 207:34]
  wire  sum_2860 = sum_2774 ^ sum_2775; // @[Mul.scala 206:34]
  wire  cout_2860 = sum_2774 & sum_2775; // @[Mul.scala 207:34]
  wire  sum_2861 = cout_2772 ^ cout_2773; // @[Mul.scala 206:34]
  wire  cout_2861 = cout_2772 & cout_2773; // @[Mul.scala 207:34]
  wire  sum_2862 = sum_2776 ^ sum_2777; // @[Mul.scala 206:34]
  wire  cout_2862 = sum_2776 & sum_2777; // @[Mul.scala 207:34]
  wire  sum_2863 = cout_2774 ^ cout_2775; // @[Mul.scala 206:34]
  wire  cout_2863 = cout_2774 & cout_2775; // @[Mul.scala 207:34]
  wire  sum_2864 = sum_2778 ^ sum_2779; // @[Mul.scala 206:34]
  wire  cout_2864 = sum_2778 & sum_2779; // @[Mul.scala 207:34]
  wire  sum_2865 = cout_2776 ^ cout_2777; // @[Mul.scala 206:34]
  wire  cout_2865 = cout_2776 & cout_2777; // @[Mul.scala 207:34]
  wire  sum_2866 = sum_2780 ^ sum_2781; // @[Mul.scala 206:34]
  wire  cout_2866 = sum_2780 & sum_2781; // @[Mul.scala 207:34]
  wire  sum_2867 = cout_2778 ^ cout_2779; // @[Mul.scala 206:34]
  wire  cout_2867 = cout_2778 & cout_2779; // @[Mul.scala 207:34]
  wire  sum_2868 = sum_2782 ^ sum_2783; // @[Mul.scala 206:34]
  wire  cout_2868 = sum_2782 & sum_2783; // @[Mul.scala 207:34]
  wire  sum_2869 = cout_2780 ^ cout_2781; // @[Mul.scala 206:34]
  wire  cout_2869 = cout_2780 & cout_2781; // @[Mul.scala 207:34]
  wire  _sum_T_3528 = sum_2784 ^ cout_2782; // @[Mul.scala 191:34]
  wire  sum_2870 = sum_2784 ^ cout_2782 ^ cout_2783; // @[Mul.scala 191:42]
  wire  cout_2870 = sum_2784 & cout_2782 | _sum_T_3528 & cout_2783; // @[Mul.scala 192:44]
  wire  sum_2871 = sum_2785 ^ cout_2784; // @[Mul.scala 206:34]
  wire  cout_2871 = sum_2785 & cout_2784; // @[Mul.scala 207:34]
  wire  sum_2872 = sum_2786 ^ cout_2785; // @[Mul.scala 206:34]
  wire  cout_2872 = sum_2786 & cout_2785; // @[Mul.scala 207:34]
  wire  sum_2873 = sum_2787 ^ cout_2786; // @[Mul.scala 206:34]
  wire  cout_2873 = sum_2787 & cout_2786; // @[Mul.scala 207:34]
  wire  sum_2874 = sum_2788 ^ cout_2787; // @[Mul.scala 206:34]
  wire  cout_2874 = sum_2788 & cout_2787; // @[Mul.scala 207:34]
  wire  sum_2875 = sum_2789 ^ cout_2788; // @[Mul.scala 206:34]
  wire  sum_2907 = sum_2821 ^ cout_2820; // @[Mul.scala 206:34]
  wire  cout_2907 = sum_2821 & cout_2820; // @[Mul.scala 207:34]
  wire  sum_2908 = sum_2822 ^ cout_2821; // @[Mul.scala 206:34]
  wire  cout_2908 = sum_2822 & cout_2821; // @[Mul.scala 207:34]
  wire  sum_2909 = sum_2823 ^ cout_2822; // @[Mul.scala 206:34]
  wire  cout_2909 = sum_2823 & cout_2822; // @[Mul.scala 207:34]
  wire  _sum_T_3569 = sum_2824 ^ sum_2825; // @[Mul.scala 191:34]
  wire  sum_2910 = sum_2824 ^ sum_2825 ^ cout_2823; // @[Mul.scala 191:42]
  wire  cout_2910 = sum_2824 & sum_2825 | _sum_T_3569 & cout_2823; // @[Mul.scala 192:44]
  wire  sum_2911 = sum_2826 ^ sum_2827; // @[Mul.scala 206:34]
  wire  cout_2911 = sum_2826 & sum_2827; // @[Mul.scala 207:34]
  wire  sum_2912 = cout_2824 ^ cout_2825; // @[Mul.scala 206:34]
  wire  cout_2912 = cout_2824 & cout_2825; // @[Mul.scala 207:34]
  wire  sum_2913 = sum_2828 ^ sum_2829; // @[Mul.scala 206:34]
  wire  cout_2913 = sum_2828 & sum_2829; // @[Mul.scala 207:34]
  wire  sum_2914 = cout_2826 ^ cout_2827; // @[Mul.scala 206:34]
  wire  cout_2914 = cout_2826 & cout_2827; // @[Mul.scala 207:34]
  wire  sum_2915 = sum_2830 ^ sum_2831; // @[Mul.scala 206:34]
  wire  cout_2915 = sum_2830 & sum_2831; // @[Mul.scala 207:34]
  wire  sum_2916 = cout_2828 ^ cout_2829; // @[Mul.scala 206:34]
  wire  cout_2916 = cout_2828 & cout_2829; // @[Mul.scala 207:34]
  wire  sum_2917 = sum_2832 ^ sum_2833; // @[Mul.scala 206:34]
  wire  cout_2917 = sum_2832 & sum_2833; // @[Mul.scala 207:34]
  wire  sum_2918 = cout_2830 ^ cout_2831; // @[Mul.scala 206:34]
  wire  cout_2918 = cout_2830 & cout_2831; // @[Mul.scala 207:34]
  wire  sum_2919 = sum_2834 ^ sum_2835; // @[Mul.scala 206:34]
  wire  cout_2919 = sum_2834 & sum_2835; // @[Mul.scala 207:34]
  wire  sum_2920 = cout_2832 ^ cout_2833; // @[Mul.scala 206:34]
  wire  cout_2920 = cout_2832 & cout_2833; // @[Mul.scala 207:34]
  wire  sum_2921 = sum_2836 ^ sum_2837; // @[Mul.scala 206:34]
  wire  cout_2921 = sum_2836 & sum_2837; // @[Mul.scala 207:34]
  wire  sum_2922 = cout_2834 ^ cout_2835; // @[Mul.scala 206:34]
  wire  cout_2922 = cout_2834 & cout_2835; // @[Mul.scala 207:34]
  wire  sum_2923 = sum_2838 ^ sum_2839; // @[Mul.scala 206:34]
  wire  cout_2923 = sum_2838 & sum_2839; // @[Mul.scala 207:34]
  wire  sum_2924 = cout_2836 ^ cout_2837; // @[Mul.scala 206:34]
  wire  cout_2924 = cout_2836 & cout_2837; // @[Mul.scala 207:34]
  wire  sum_2925 = sum_2840 ^ sum_2841; // @[Mul.scala 206:34]
  wire  cout_2925 = sum_2840 & sum_2841; // @[Mul.scala 207:34]
  wire  sum_2926 = cout_2838 ^ cout_2839; // @[Mul.scala 206:34]
  wire  cout_2926 = cout_2838 & cout_2839; // @[Mul.scala 207:34]
  wire  sum_2927 = sum_2842 ^ sum_2843; // @[Mul.scala 206:34]
  wire  cout_2927 = sum_2842 & sum_2843; // @[Mul.scala 207:34]
  wire  sum_2928 = cout_2840 ^ cout_2841; // @[Mul.scala 206:34]
  wire  cout_2928 = cout_2840 & cout_2841; // @[Mul.scala 207:34]
  wire  sum_2929 = sum_2844 ^ sum_2845; // @[Mul.scala 206:34]
  wire  cout_2929 = sum_2844 & sum_2845; // @[Mul.scala 207:34]
  wire  sum_2930 = cout_2842 ^ cout_2843; // @[Mul.scala 206:34]
  wire  cout_2930 = cout_2842 & cout_2843; // @[Mul.scala 207:34]
  wire  sum_2931 = sum_2846 ^ sum_2847; // @[Mul.scala 206:34]
  wire  cout_2931 = sum_2846 & sum_2847; // @[Mul.scala 207:34]
  wire  sum_2932 = cout_2844 ^ cout_2845; // @[Mul.scala 206:34]
  wire  cout_2932 = cout_2844 & cout_2845; // @[Mul.scala 207:34]
  wire  sum_2933 = sum_2848 ^ sum_2849; // @[Mul.scala 206:34]
  wire  cout_2933 = sum_2848 & sum_2849; // @[Mul.scala 207:34]
  wire  sum_2934 = cout_2846 ^ cout_2847; // @[Mul.scala 206:34]
  wire  cout_2934 = cout_2846 & cout_2847; // @[Mul.scala 207:34]
  wire  sum_2935 = sum_2850 ^ sum_2851; // @[Mul.scala 206:34]
  wire  cout_2935 = sum_2850 & sum_2851; // @[Mul.scala 207:34]
  wire  sum_2936 = cout_2848 ^ cout_2849; // @[Mul.scala 206:34]
  wire  cout_2936 = cout_2848 & cout_2849; // @[Mul.scala 207:34]
  wire  sum_2937 = sum_2852 ^ sum_2853; // @[Mul.scala 206:34]
  wire  cout_2937 = sum_2852 & sum_2853; // @[Mul.scala 207:34]
  wire  sum_2938 = cout_2850 ^ cout_2851; // @[Mul.scala 206:34]
  wire  cout_2938 = cout_2850 & cout_2851; // @[Mul.scala 207:34]
  wire  sum_2939 = sum_2854 ^ sum_2855; // @[Mul.scala 206:34]
  wire  cout_2939 = sum_2854 & sum_2855; // @[Mul.scala 207:34]
  wire  sum_2940 = cout_2852 ^ cout_2853; // @[Mul.scala 206:34]
  wire  cout_2940 = cout_2852 & cout_2853; // @[Mul.scala 207:34]
  wire  sum_2941 = sum_2856 ^ sum_2857; // @[Mul.scala 206:34]
  wire  cout_2941 = sum_2856 & sum_2857; // @[Mul.scala 207:34]
  wire  sum_2942 = cout_2854 ^ cout_2855; // @[Mul.scala 206:34]
  wire  cout_2942 = cout_2854 & cout_2855; // @[Mul.scala 207:34]
  wire  sum_2943 = sum_2858 ^ sum_2859; // @[Mul.scala 206:34]
  wire  cout_2943 = sum_2858 & sum_2859; // @[Mul.scala 207:34]
  wire  sum_2944 = cout_2856 ^ cout_2857; // @[Mul.scala 206:34]
  wire  cout_2944 = cout_2856 & cout_2857; // @[Mul.scala 207:34]
  wire  sum_2945 = sum_2860 ^ sum_2861; // @[Mul.scala 206:34]
  wire  cout_2945 = sum_2860 & sum_2861; // @[Mul.scala 207:34]
  wire  sum_2946 = cout_2858 ^ cout_2859; // @[Mul.scala 206:34]
  wire  cout_2946 = cout_2858 & cout_2859; // @[Mul.scala 207:34]
  wire  sum_2947 = sum_2862 ^ sum_2863; // @[Mul.scala 206:34]
  wire  cout_2947 = sum_2862 & sum_2863; // @[Mul.scala 207:34]
  wire  sum_2948 = cout_2860 ^ cout_2861; // @[Mul.scala 206:34]
  wire  cout_2948 = cout_2860 & cout_2861; // @[Mul.scala 207:34]
  wire  sum_2949 = sum_2864 ^ sum_2865; // @[Mul.scala 206:34]
  wire  cout_2949 = sum_2864 & sum_2865; // @[Mul.scala 207:34]
  wire  sum_2950 = cout_2862 ^ cout_2863; // @[Mul.scala 206:34]
  wire  cout_2950 = cout_2862 & cout_2863; // @[Mul.scala 207:34]
  wire  sum_2951 = sum_2866 ^ sum_2867; // @[Mul.scala 206:34]
  wire  cout_2951 = sum_2866 & sum_2867; // @[Mul.scala 207:34]
  wire  sum_2952 = cout_2864 ^ cout_2865; // @[Mul.scala 206:34]
  wire  cout_2952 = cout_2864 & cout_2865; // @[Mul.scala 207:34]
  wire  sum_2953 = sum_2868 ^ sum_2869; // @[Mul.scala 206:34]
  wire  cout_2953 = sum_2868 & sum_2869; // @[Mul.scala 207:34]
  wire  sum_2954 = cout_2866 ^ cout_2867; // @[Mul.scala 206:34]
  wire  cout_2954 = cout_2866 & cout_2867; // @[Mul.scala 207:34]
  wire  _sum_T_3615 = sum_2870 ^ cout_2868; // @[Mul.scala 191:34]
  wire  sum_2955 = sum_2870 ^ cout_2868 ^ cout_2869; // @[Mul.scala 191:42]
  wire  cout_2955 = sum_2870 & cout_2868 | _sum_T_3615 & cout_2869; // @[Mul.scala 192:44]
  wire  sum_2956 = sum_2871 ^ cout_2870; // @[Mul.scala 206:34]
  wire  cout_2956 = sum_2871 & cout_2870; // @[Mul.scala 207:34]
  wire  sum_2957 = sum_2872 ^ cout_2871; // @[Mul.scala 206:34]
  wire  cout_2957 = sum_2872 & cout_2871; // @[Mul.scala 207:34]
  wire  sum_2958 = sum_2873 ^ cout_2872; // @[Mul.scala 206:34]
  wire  cout_2958 = sum_2873 & cout_2872; // @[Mul.scala 207:34]
  wire  sum_2959 = sum_2874 ^ cout_2873; // @[Mul.scala 206:34]
  wire  cout_2959 = sum_2874 & cout_2873; // @[Mul.scala 207:34]
  wire  sum_2960 = sum_2875 ^ cout_2874; // @[Mul.scala 206:34]
  wire  sum_2993 = sum_2908 ^ cout_2907; // @[Mul.scala 206:34]
  wire  cout_2993 = sum_2908 & cout_2907; // @[Mul.scala 207:34]
  wire  sum_2994 = sum_2909 ^ cout_2908; // @[Mul.scala 206:34]
  wire  cout_2994 = sum_2909 & cout_2908; // @[Mul.scala 207:34]
  wire  sum_2995 = sum_2910 ^ cout_2909; // @[Mul.scala 206:34]
  wire  cout_2995 = sum_2910 & cout_2909; // @[Mul.scala 207:34]
  wire  _sum_T_3657 = sum_2911 ^ sum_2912; // @[Mul.scala 191:34]
  wire  sum_2996 = sum_2911 ^ sum_2912 ^ cout_2910; // @[Mul.scala 191:42]
  wire  cout_2996 = sum_2911 & sum_2912 | _sum_T_3657 & cout_2910; // @[Mul.scala 192:44]
  wire  sum_2997 = sum_2913 ^ sum_2914; // @[Mul.scala 206:34]
  wire  cout_2997 = sum_2913 & sum_2914; // @[Mul.scala 207:34]
  wire  sum_2998 = cout_2911 ^ cout_2912; // @[Mul.scala 206:34]
  wire  cout_2998 = cout_2911 & cout_2912; // @[Mul.scala 207:34]
  wire  sum_2999 = sum_2915 ^ sum_2916; // @[Mul.scala 206:34]
  wire  cout_2999 = sum_2915 & sum_2916; // @[Mul.scala 207:34]
  wire  sum_3000 = cout_2913 ^ cout_2914; // @[Mul.scala 206:34]
  wire  cout_3000 = cout_2913 & cout_2914; // @[Mul.scala 207:34]
  wire  sum_3001 = sum_2917 ^ sum_2918; // @[Mul.scala 206:34]
  wire  cout_3001 = sum_2917 & sum_2918; // @[Mul.scala 207:34]
  wire  sum_3002 = cout_2915 ^ cout_2916; // @[Mul.scala 206:34]
  wire  cout_3002 = cout_2915 & cout_2916; // @[Mul.scala 207:34]
  wire  sum_3003 = sum_2919 ^ sum_2920; // @[Mul.scala 206:34]
  wire  cout_3003 = sum_2919 & sum_2920; // @[Mul.scala 207:34]
  wire  sum_3004 = cout_2917 ^ cout_2918; // @[Mul.scala 206:34]
  wire  cout_3004 = cout_2917 & cout_2918; // @[Mul.scala 207:34]
  wire  sum_3005 = sum_2921 ^ sum_2922; // @[Mul.scala 206:34]
  wire  cout_3005 = sum_2921 & sum_2922; // @[Mul.scala 207:34]
  wire  sum_3006 = cout_2919 ^ cout_2920; // @[Mul.scala 206:34]
  wire  cout_3006 = cout_2919 & cout_2920; // @[Mul.scala 207:34]
  wire  sum_3007 = sum_2923 ^ sum_2924; // @[Mul.scala 206:34]
  wire  cout_3007 = sum_2923 & sum_2924; // @[Mul.scala 207:34]
  wire  sum_3008 = cout_2921 ^ cout_2922; // @[Mul.scala 206:34]
  wire  cout_3008 = cout_2921 & cout_2922; // @[Mul.scala 207:34]
  wire  sum_3009 = sum_2925 ^ sum_2926; // @[Mul.scala 206:34]
  wire  cout_3009 = sum_2925 & sum_2926; // @[Mul.scala 207:34]
  wire  sum_3010 = cout_2923 ^ cout_2924; // @[Mul.scala 206:34]
  wire  cout_3010 = cout_2923 & cout_2924; // @[Mul.scala 207:34]
  wire  sum_3011 = sum_2927 ^ sum_2928; // @[Mul.scala 206:34]
  wire  cout_3011 = sum_2927 & sum_2928; // @[Mul.scala 207:34]
  wire  sum_3012 = cout_2925 ^ cout_2926; // @[Mul.scala 206:34]
  wire  cout_3012 = cout_2925 & cout_2926; // @[Mul.scala 207:34]
  wire  sum_3013 = sum_2929 ^ sum_2930; // @[Mul.scala 206:34]
  wire  cout_3013 = sum_2929 & sum_2930; // @[Mul.scala 207:34]
  wire  sum_3014 = cout_2927 ^ cout_2928; // @[Mul.scala 206:34]
  wire  cout_3014 = cout_2927 & cout_2928; // @[Mul.scala 207:34]
  wire  sum_3015 = sum_2931 ^ sum_2932; // @[Mul.scala 206:34]
  wire  cout_3015 = sum_2931 & sum_2932; // @[Mul.scala 207:34]
  wire  sum_3016 = cout_2929 ^ cout_2930; // @[Mul.scala 206:34]
  wire  cout_3016 = cout_2929 & cout_2930; // @[Mul.scala 207:34]
  wire  sum_3017 = sum_2933 ^ sum_2934; // @[Mul.scala 206:34]
  wire  cout_3017 = sum_2933 & sum_2934; // @[Mul.scala 207:34]
  wire  sum_3018 = cout_2931 ^ cout_2932; // @[Mul.scala 206:34]
  wire  cout_3018 = cout_2931 & cout_2932; // @[Mul.scala 207:34]
  wire  sum_3019 = sum_2935 ^ sum_2936; // @[Mul.scala 206:34]
  wire  cout_3019 = sum_2935 & sum_2936; // @[Mul.scala 207:34]
  wire  sum_3020 = cout_2933 ^ cout_2934; // @[Mul.scala 206:34]
  wire  cout_3020 = cout_2933 & cout_2934; // @[Mul.scala 207:34]
  wire  sum_3021 = sum_2937 ^ sum_2938; // @[Mul.scala 206:34]
  wire  cout_3021 = sum_2937 & sum_2938; // @[Mul.scala 207:34]
  wire  sum_3022 = cout_2935 ^ cout_2936; // @[Mul.scala 206:34]
  wire  cout_3022 = cout_2935 & cout_2936; // @[Mul.scala 207:34]
  wire  sum_3023 = sum_2939 ^ sum_2940; // @[Mul.scala 206:34]
  wire  cout_3023 = sum_2939 & sum_2940; // @[Mul.scala 207:34]
  wire  sum_3024 = cout_2937 ^ cout_2938; // @[Mul.scala 206:34]
  wire  cout_3024 = cout_2937 & cout_2938; // @[Mul.scala 207:34]
  wire  sum_3025 = sum_2941 ^ sum_2942; // @[Mul.scala 206:34]
  wire  cout_3025 = sum_2941 & sum_2942; // @[Mul.scala 207:34]
  wire  sum_3026 = cout_2939 ^ cout_2940; // @[Mul.scala 206:34]
  wire  cout_3026 = cout_2939 & cout_2940; // @[Mul.scala 207:34]
  wire  sum_3027 = sum_2943 ^ sum_2944; // @[Mul.scala 206:34]
  wire  cout_3027 = sum_2943 & sum_2944; // @[Mul.scala 207:34]
  wire  sum_3028 = cout_2941 ^ cout_2942; // @[Mul.scala 206:34]
  wire  cout_3028 = cout_2941 & cout_2942; // @[Mul.scala 207:34]
  wire  sum_3029 = sum_2945 ^ sum_2946; // @[Mul.scala 206:34]
  wire  cout_3029 = sum_2945 & sum_2946; // @[Mul.scala 207:34]
  wire  sum_3030 = cout_2943 ^ cout_2944; // @[Mul.scala 206:34]
  wire  cout_3030 = cout_2943 & cout_2944; // @[Mul.scala 207:34]
  wire  sum_3031 = sum_2947 ^ sum_2948; // @[Mul.scala 206:34]
  wire  cout_3031 = sum_2947 & sum_2948; // @[Mul.scala 207:34]
  wire  sum_3032 = cout_2945 ^ cout_2946; // @[Mul.scala 206:34]
  wire  cout_3032 = cout_2945 & cout_2946; // @[Mul.scala 207:34]
  wire  sum_3033 = sum_2949 ^ sum_2950; // @[Mul.scala 206:34]
  wire  cout_3033 = sum_2949 & sum_2950; // @[Mul.scala 207:34]
  wire  sum_3034 = cout_2947 ^ cout_2948; // @[Mul.scala 206:34]
  wire  cout_3034 = cout_2947 & cout_2948; // @[Mul.scala 207:34]
  wire  sum_3035 = sum_2951 ^ sum_2952; // @[Mul.scala 206:34]
  wire  cout_3035 = sum_2951 & sum_2952; // @[Mul.scala 207:34]
  wire  sum_3036 = cout_2949 ^ cout_2950; // @[Mul.scala 206:34]
  wire  cout_3036 = cout_2949 & cout_2950; // @[Mul.scala 207:34]
  wire  sum_3037 = sum_2953 ^ sum_2954; // @[Mul.scala 206:34]
  wire  cout_3037 = sum_2953 & sum_2954; // @[Mul.scala 207:34]
  wire  sum_3038 = cout_2951 ^ cout_2952; // @[Mul.scala 206:34]
  wire  cout_3038 = cout_2951 & cout_2952; // @[Mul.scala 207:34]
  wire  _sum_T_3701 = sum_2955 ^ cout_2953; // @[Mul.scala 191:34]
  wire  sum_3039 = sum_2955 ^ cout_2953 ^ cout_2954; // @[Mul.scala 191:42]
  wire  cout_3039 = sum_2955 & cout_2953 | _sum_T_3701 & cout_2954; // @[Mul.scala 192:44]
  wire  sum_3040 = sum_2956 ^ cout_2955; // @[Mul.scala 206:34]
  wire  cout_3040 = sum_2956 & cout_2955; // @[Mul.scala 207:34]
  wire  sum_3041 = sum_2957 ^ cout_2956; // @[Mul.scala 206:34]
  wire  cout_3041 = sum_2957 & cout_2956; // @[Mul.scala 207:34]
  wire  sum_3042 = sum_2958 ^ cout_2957; // @[Mul.scala 206:34]
  wire  cout_3042 = sum_2958 & cout_2957; // @[Mul.scala 207:34]
  wire  sum_3043 = sum_2959 ^ cout_2958; // @[Mul.scala 206:34]
  wire  cout_3043 = sum_2959 & cout_2958; // @[Mul.scala 207:34]
  wire  sum_3044 = sum_2960 ^ cout_2959; // @[Mul.scala 206:34]
  wire  sum_3078 = sum_2994 ^ cout_2993; // @[Mul.scala 206:34]
  wire  cout_3078 = sum_2994 & cout_2993; // @[Mul.scala 207:34]
  wire  sum_3079 = sum_2995 ^ cout_2994; // @[Mul.scala 206:34]
  wire  cout_3079 = sum_2995 & cout_2994; // @[Mul.scala 207:34]
  wire  sum_3080 = sum_2996 ^ cout_2995; // @[Mul.scala 206:34]
  wire  cout_3080 = sum_2996 & cout_2995; // @[Mul.scala 207:34]
  wire  _sum_T_3744 = sum_2997 ^ sum_2998; // @[Mul.scala 191:34]
  wire  sum_3081 = sum_2997 ^ sum_2998 ^ cout_2996; // @[Mul.scala 191:42]
  wire  cout_3081 = sum_2997 & sum_2998 | _sum_T_3744 & cout_2996; // @[Mul.scala 192:44]
  wire  sum_3082 = sum_2999 ^ sum_3000; // @[Mul.scala 206:34]
  wire  cout_3082 = sum_2999 & sum_3000; // @[Mul.scala 207:34]
  wire  sum_3083 = cout_2997 ^ cout_2998; // @[Mul.scala 206:34]
  wire  cout_3083 = cout_2997 & cout_2998; // @[Mul.scala 207:34]
  wire  sum_3084 = sum_3001 ^ sum_3002; // @[Mul.scala 206:34]
  wire  cout_3084 = sum_3001 & sum_3002; // @[Mul.scala 207:34]
  wire  sum_3085 = cout_2999 ^ cout_3000; // @[Mul.scala 206:34]
  wire  cout_3085 = cout_2999 & cout_3000; // @[Mul.scala 207:34]
  wire  sum_3086 = sum_3003 ^ sum_3004; // @[Mul.scala 206:34]
  wire  cout_3086 = sum_3003 & sum_3004; // @[Mul.scala 207:34]
  wire  sum_3087 = cout_3001 ^ cout_3002; // @[Mul.scala 206:34]
  wire  cout_3087 = cout_3001 & cout_3002; // @[Mul.scala 207:34]
  wire  sum_3088 = sum_3005 ^ sum_3006; // @[Mul.scala 206:34]
  wire  cout_3088 = sum_3005 & sum_3006; // @[Mul.scala 207:34]
  wire  sum_3089 = cout_3003 ^ cout_3004; // @[Mul.scala 206:34]
  wire  cout_3089 = cout_3003 & cout_3004; // @[Mul.scala 207:34]
  wire  sum_3090 = sum_3007 ^ sum_3008; // @[Mul.scala 206:34]
  wire  cout_3090 = sum_3007 & sum_3008; // @[Mul.scala 207:34]
  wire  sum_3091 = cout_3005 ^ cout_3006; // @[Mul.scala 206:34]
  wire  cout_3091 = cout_3005 & cout_3006; // @[Mul.scala 207:34]
  wire  sum_3092 = sum_3009 ^ sum_3010; // @[Mul.scala 206:34]
  wire  cout_3092 = sum_3009 & sum_3010; // @[Mul.scala 207:34]
  wire  sum_3093 = cout_3007 ^ cout_3008; // @[Mul.scala 206:34]
  wire  cout_3093 = cout_3007 & cout_3008; // @[Mul.scala 207:34]
  wire  sum_3094 = sum_3011 ^ sum_3012; // @[Mul.scala 206:34]
  wire  cout_3094 = sum_3011 & sum_3012; // @[Mul.scala 207:34]
  wire  sum_3095 = cout_3009 ^ cout_3010; // @[Mul.scala 206:34]
  wire  cout_3095 = cout_3009 & cout_3010; // @[Mul.scala 207:34]
  wire  sum_3096 = sum_3013 ^ sum_3014; // @[Mul.scala 206:34]
  wire  cout_3096 = sum_3013 & sum_3014; // @[Mul.scala 207:34]
  wire  sum_3097 = cout_3011 ^ cout_3012; // @[Mul.scala 206:34]
  wire  cout_3097 = cout_3011 & cout_3012; // @[Mul.scala 207:34]
  wire  sum_3098 = sum_3015 ^ sum_3016; // @[Mul.scala 206:34]
  wire  cout_3098 = sum_3015 & sum_3016; // @[Mul.scala 207:34]
  wire  sum_3099 = cout_3013 ^ cout_3014; // @[Mul.scala 206:34]
  wire  cout_3099 = cout_3013 & cout_3014; // @[Mul.scala 207:34]
  wire  sum_3100 = sum_3017 ^ sum_3018; // @[Mul.scala 206:34]
  wire  cout_3100 = sum_3017 & sum_3018; // @[Mul.scala 207:34]
  wire  sum_3101 = cout_3015 ^ cout_3016; // @[Mul.scala 206:34]
  wire  cout_3101 = cout_3015 & cout_3016; // @[Mul.scala 207:34]
  wire  sum_3102 = sum_3019 ^ sum_3020; // @[Mul.scala 206:34]
  wire  cout_3102 = sum_3019 & sum_3020; // @[Mul.scala 207:34]
  wire  sum_3103 = cout_3017 ^ cout_3018; // @[Mul.scala 206:34]
  wire  cout_3103 = cout_3017 & cout_3018; // @[Mul.scala 207:34]
  wire  sum_3104 = sum_3021 ^ sum_3022; // @[Mul.scala 206:34]
  wire  cout_3104 = sum_3021 & sum_3022; // @[Mul.scala 207:34]
  wire  sum_3105 = cout_3019 ^ cout_3020; // @[Mul.scala 206:34]
  wire  cout_3105 = cout_3019 & cout_3020; // @[Mul.scala 207:34]
  wire  sum_3106 = sum_3023 ^ sum_3024; // @[Mul.scala 206:34]
  wire  cout_3106 = sum_3023 & sum_3024; // @[Mul.scala 207:34]
  wire  sum_3107 = cout_3021 ^ cout_3022; // @[Mul.scala 206:34]
  wire  cout_3107 = cout_3021 & cout_3022; // @[Mul.scala 207:34]
  wire  sum_3108 = sum_3025 ^ sum_3026; // @[Mul.scala 206:34]
  wire  cout_3108 = sum_3025 & sum_3026; // @[Mul.scala 207:34]
  wire  sum_3109 = cout_3023 ^ cout_3024; // @[Mul.scala 206:34]
  wire  cout_3109 = cout_3023 & cout_3024; // @[Mul.scala 207:34]
  wire  sum_3110 = sum_3027 ^ sum_3028; // @[Mul.scala 206:34]
  wire  cout_3110 = sum_3027 & sum_3028; // @[Mul.scala 207:34]
  wire  sum_3111 = cout_3025 ^ cout_3026; // @[Mul.scala 206:34]
  wire  cout_3111 = cout_3025 & cout_3026; // @[Mul.scala 207:34]
  wire  sum_3112 = sum_3029 ^ sum_3030; // @[Mul.scala 206:34]
  wire  cout_3112 = sum_3029 & sum_3030; // @[Mul.scala 207:34]
  wire  sum_3113 = cout_3027 ^ cout_3028; // @[Mul.scala 206:34]
  wire  cout_3113 = cout_3027 & cout_3028; // @[Mul.scala 207:34]
  wire  sum_3114 = sum_3031 ^ sum_3032; // @[Mul.scala 206:34]
  wire  cout_3114 = sum_3031 & sum_3032; // @[Mul.scala 207:34]
  wire  sum_3115 = cout_3029 ^ cout_3030; // @[Mul.scala 206:34]
  wire  cout_3115 = cout_3029 & cout_3030; // @[Mul.scala 207:34]
  wire  sum_3116 = sum_3033 ^ sum_3034; // @[Mul.scala 206:34]
  wire  cout_3116 = sum_3033 & sum_3034; // @[Mul.scala 207:34]
  wire  sum_3117 = cout_3031 ^ cout_3032; // @[Mul.scala 206:34]
  wire  cout_3117 = cout_3031 & cout_3032; // @[Mul.scala 207:34]
  wire  sum_3118 = sum_3035 ^ sum_3036; // @[Mul.scala 206:34]
  wire  cout_3118 = sum_3035 & sum_3036; // @[Mul.scala 207:34]
  wire  sum_3119 = cout_3033 ^ cout_3034; // @[Mul.scala 206:34]
  wire  cout_3119 = cout_3033 & cout_3034; // @[Mul.scala 207:34]
  wire  sum_3120 = sum_3037 ^ sum_3038; // @[Mul.scala 206:34]
  wire  cout_3120 = sum_3037 & sum_3038; // @[Mul.scala 207:34]
  wire  sum_3121 = cout_3035 ^ cout_3036; // @[Mul.scala 206:34]
  wire  cout_3121 = cout_3035 & cout_3036; // @[Mul.scala 207:34]
  wire  _sum_T_3786 = sum_3039 ^ cout_3037; // @[Mul.scala 191:34]
  wire  sum_3122 = sum_3039 ^ cout_3037 ^ cout_3038; // @[Mul.scala 191:42]
  wire  cout_3122 = sum_3039 & cout_3037 | _sum_T_3786 & cout_3038; // @[Mul.scala 192:44]
  wire  sum_3123 = sum_3040 ^ cout_3039; // @[Mul.scala 206:34]
  wire  cout_3123 = sum_3040 & cout_3039; // @[Mul.scala 207:34]
  wire  sum_3124 = sum_3041 ^ cout_3040; // @[Mul.scala 206:34]
  wire  cout_3124 = sum_3041 & cout_3040; // @[Mul.scala 207:34]
  wire  sum_3125 = sum_3042 ^ cout_3041; // @[Mul.scala 206:34]
  wire  cout_3125 = sum_3042 & cout_3041; // @[Mul.scala 207:34]
  wire  sum_3126 = sum_3043 ^ cout_3042; // @[Mul.scala 206:34]
  wire  cout_3126 = sum_3043 & cout_3042; // @[Mul.scala 207:34]
  wire  sum_3127 = sum_3044 ^ cout_3043; // @[Mul.scala 206:34]
  wire  sum_3162 = sum_3079 ^ cout_3078; // @[Mul.scala 206:34]
  wire  cout_3162 = sum_3079 & cout_3078; // @[Mul.scala 207:34]
  wire  sum_3163 = sum_3080 ^ cout_3079; // @[Mul.scala 206:34]
  wire  cout_3163 = sum_3080 & cout_3079; // @[Mul.scala 207:34]
  wire  sum_3164 = sum_3081 ^ cout_3080; // @[Mul.scala 206:34]
  wire  cout_3164 = sum_3081 & cout_3080; // @[Mul.scala 207:34]
  wire  _sum_T_3830 = sum_3082 ^ sum_3083; // @[Mul.scala 191:34]
  wire  sum_3165 = sum_3082 ^ sum_3083 ^ cout_3081; // @[Mul.scala 191:42]
  wire  cout_3165 = sum_3082 & sum_3083 | _sum_T_3830 & cout_3081; // @[Mul.scala 192:44]
  wire  sum_3166 = sum_3084 ^ sum_3085; // @[Mul.scala 206:34]
  wire  cout_3166 = sum_3084 & sum_3085; // @[Mul.scala 207:34]
  wire  sum_3167 = cout_3082 ^ cout_3083; // @[Mul.scala 206:34]
  wire  cout_3167 = cout_3082 & cout_3083; // @[Mul.scala 207:34]
  wire  sum_3168 = sum_3086 ^ sum_3087; // @[Mul.scala 206:34]
  wire  cout_3168 = sum_3086 & sum_3087; // @[Mul.scala 207:34]
  wire  sum_3169 = cout_3084 ^ cout_3085; // @[Mul.scala 206:34]
  wire  cout_3169 = cout_3084 & cout_3085; // @[Mul.scala 207:34]
  wire  sum_3170 = sum_3088 ^ sum_3089; // @[Mul.scala 206:34]
  wire  cout_3170 = sum_3088 & sum_3089; // @[Mul.scala 207:34]
  wire  sum_3171 = cout_3086 ^ cout_3087; // @[Mul.scala 206:34]
  wire  cout_3171 = cout_3086 & cout_3087; // @[Mul.scala 207:34]
  wire  sum_3172 = sum_3090 ^ sum_3091; // @[Mul.scala 206:34]
  wire  cout_3172 = sum_3090 & sum_3091; // @[Mul.scala 207:34]
  wire  sum_3173 = cout_3088 ^ cout_3089; // @[Mul.scala 206:34]
  wire  cout_3173 = cout_3088 & cout_3089; // @[Mul.scala 207:34]
  wire  sum_3174 = sum_3092 ^ sum_3093; // @[Mul.scala 206:34]
  wire  cout_3174 = sum_3092 & sum_3093; // @[Mul.scala 207:34]
  wire  sum_3175 = cout_3090 ^ cout_3091; // @[Mul.scala 206:34]
  wire  cout_3175 = cout_3090 & cout_3091; // @[Mul.scala 207:34]
  wire  sum_3176 = sum_3094 ^ sum_3095; // @[Mul.scala 206:34]
  wire  cout_3176 = sum_3094 & sum_3095; // @[Mul.scala 207:34]
  wire  sum_3177 = cout_3092 ^ cout_3093; // @[Mul.scala 206:34]
  wire  cout_3177 = cout_3092 & cout_3093; // @[Mul.scala 207:34]
  wire  sum_3178 = sum_3096 ^ sum_3097; // @[Mul.scala 206:34]
  wire  cout_3178 = sum_3096 & sum_3097; // @[Mul.scala 207:34]
  wire  sum_3179 = cout_3094 ^ cout_3095; // @[Mul.scala 206:34]
  wire  cout_3179 = cout_3094 & cout_3095; // @[Mul.scala 207:34]
  wire  sum_3180 = sum_3098 ^ sum_3099; // @[Mul.scala 206:34]
  wire  cout_3180 = sum_3098 & sum_3099; // @[Mul.scala 207:34]
  wire  sum_3181 = cout_3096 ^ cout_3097; // @[Mul.scala 206:34]
  wire  cout_3181 = cout_3096 & cout_3097; // @[Mul.scala 207:34]
  wire  sum_3182 = sum_3100 ^ sum_3101; // @[Mul.scala 206:34]
  wire  cout_3182 = sum_3100 & sum_3101; // @[Mul.scala 207:34]
  wire  sum_3183 = cout_3098 ^ cout_3099; // @[Mul.scala 206:34]
  wire  cout_3183 = cout_3098 & cout_3099; // @[Mul.scala 207:34]
  wire  sum_3184 = sum_3102 ^ sum_3103; // @[Mul.scala 206:34]
  wire  cout_3184 = sum_3102 & sum_3103; // @[Mul.scala 207:34]
  wire  sum_3185 = cout_3100 ^ cout_3101; // @[Mul.scala 206:34]
  wire  cout_3185 = cout_3100 & cout_3101; // @[Mul.scala 207:34]
  wire  sum_3186 = sum_3104 ^ sum_3105; // @[Mul.scala 206:34]
  wire  cout_3186 = sum_3104 & sum_3105; // @[Mul.scala 207:34]
  wire  sum_3187 = cout_3102 ^ cout_3103; // @[Mul.scala 206:34]
  wire  cout_3187 = cout_3102 & cout_3103; // @[Mul.scala 207:34]
  wire  sum_3188 = sum_3106 ^ sum_3107; // @[Mul.scala 206:34]
  wire  cout_3188 = sum_3106 & sum_3107; // @[Mul.scala 207:34]
  wire  sum_3189 = cout_3104 ^ cout_3105; // @[Mul.scala 206:34]
  wire  cout_3189 = cout_3104 & cout_3105; // @[Mul.scala 207:34]
  wire  sum_3190 = sum_3108 ^ sum_3109; // @[Mul.scala 206:34]
  wire  cout_3190 = sum_3108 & sum_3109; // @[Mul.scala 207:34]
  wire  sum_3191 = cout_3106 ^ cout_3107; // @[Mul.scala 206:34]
  wire  cout_3191 = cout_3106 & cout_3107; // @[Mul.scala 207:34]
  wire  sum_3192 = sum_3110 ^ sum_3111; // @[Mul.scala 206:34]
  wire  cout_3192 = sum_3110 & sum_3111; // @[Mul.scala 207:34]
  wire  sum_3193 = cout_3108 ^ cout_3109; // @[Mul.scala 206:34]
  wire  cout_3193 = cout_3108 & cout_3109; // @[Mul.scala 207:34]
  wire  sum_3194 = sum_3112 ^ sum_3113; // @[Mul.scala 206:34]
  wire  cout_3194 = sum_3112 & sum_3113; // @[Mul.scala 207:34]
  wire  sum_3195 = cout_3110 ^ cout_3111; // @[Mul.scala 206:34]
  wire  cout_3195 = cout_3110 & cout_3111; // @[Mul.scala 207:34]
  wire  sum_3196 = sum_3114 ^ sum_3115; // @[Mul.scala 206:34]
  wire  cout_3196 = sum_3114 & sum_3115; // @[Mul.scala 207:34]
  wire  sum_3197 = cout_3112 ^ cout_3113; // @[Mul.scala 206:34]
  wire  cout_3197 = cout_3112 & cout_3113; // @[Mul.scala 207:34]
  wire  sum_3198 = sum_3116 ^ sum_3117; // @[Mul.scala 206:34]
  wire  cout_3198 = sum_3116 & sum_3117; // @[Mul.scala 207:34]
  wire  sum_3199 = cout_3114 ^ cout_3115; // @[Mul.scala 206:34]
  wire  cout_3199 = cout_3114 & cout_3115; // @[Mul.scala 207:34]
  wire  sum_3200 = sum_3118 ^ sum_3119; // @[Mul.scala 206:34]
  wire  cout_3200 = sum_3118 & sum_3119; // @[Mul.scala 207:34]
  wire  sum_3201 = cout_3116 ^ cout_3117; // @[Mul.scala 206:34]
  wire  cout_3201 = cout_3116 & cout_3117; // @[Mul.scala 207:34]
  wire  sum_3202 = sum_3120 ^ sum_3121; // @[Mul.scala 206:34]
  wire  cout_3202 = sum_3120 & sum_3121; // @[Mul.scala 207:34]
  wire  sum_3203 = cout_3118 ^ cout_3119; // @[Mul.scala 206:34]
  wire  cout_3203 = cout_3118 & cout_3119; // @[Mul.scala 207:34]
  wire  _sum_T_3870 = sum_3122 ^ cout_3120; // @[Mul.scala 191:34]
  wire  sum_3204 = sum_3122 ^ cout_3120 ^ cout_3121; // @[Mul.scala 191:42]
  wire  cout_3204 = sum_3122 & cout_3120 | _sum_T_3870 & cout_3121; // @[Mul.scala 192:44]
  wire  sum_3205 = sum_3123 ^ cout_3122; // @[Mul.scala 206:34]
  wire  cout_3205 = sum_3123 & cout_3122; // @[Mul.scala 207:34]
  wire  sum_3206 = sum_3124 ^ cout_3123; // @[Mul.scala 206:34]
  wire  cout_3206 = sum_3124 & cout_3123; // @[Mul.scala 207:34]
  wire  sum_3207 = sum_3125 ^ cout_3124; // @[Mul.scala 206:34]
  wire  cout_3207 = sum_3125 & cout_3124; // @[Mul.scala 207:34]
  wire  sum_3208 = sum_3126 ^ cout_3125; // @[Mul.scala 206:34]
  wire  cout_3208 = sum_3126 & cout_3125; // @[Mul.scala 207:34]
  wire  sum_3209 = sum_3127 ^ cout_3126; // @[Mul.scala 206:34]
  wire  sum_3245 = sum_3163 ^ cout_3162; // @[Mul.scala 206:34]
  wire  cout_3245 = sum_3163 & cout_3162; // @[Mul.scala 207:34]
  wire  sum_3246 = sum_3164 ^ cout_3163; // @[Mul.scala 206:34]
  wire  cout_3246 = sum_3164 & cout_3163; // @[Mul.scala 207:34]
  wire  sum_3247 = sum_3165 ^ cout_3164; // @[Mul.scala 206:34]
  wire  cout_3247 = sum_3165 & cout_3164; // @[Mul.scala 207:34]
  wire  _sum_T_3915 = sum_3166 ^ sum_3167; // @[Mul.scala 191:34]
  wire  sum_3248 = sum_3166 ^ sum_3167 ^ cout_3165; // @[Mul.scala 191:42]
  wire  cout_3248 = sum_3166 & sum_3167 | _sum_T_3915 & cout_3165; // @[Mul.scala 192:44]
  wire  sum_3249 = sum_3168 ^ sum_3169; // @[Mul.scala 206:34]
  wire  cout_3249 = sum_3168 & sum_3169; // @[Mul.scala 207:34]
  wire  sum_3250 = cout_3166 ^ cout_3167; // @[Mul.scala 206:34]
  wire  cout_3250 = cout_3166 & cout_3167; // @[Mul.scala 207:34]
  wire  sum_3251 = sum_3170 ^ sum_3171; // @[Mul.scala 206:34]
  wire  cout_3251 = sum_3170 & sum_3171; // @[Mul.scala 207:34]
  wire  sum_3252 = cout_3168 ^ cout_3169; // @[Mul.scala 206:34]
  wire  cout_3252 = cout_3168 & cout_3169; // @[Mul.scala 207:34]
  wire  sum_3253 = sum_3172 ^ sum_3173; // @[Mul.scala 206:34]
  wire  cout_3253 = sum_3172 & sum_3173; // @[Mul.scala 207:34]
  wire  sum_3254 = cout_3170 ^ cout_3171; // @[Mul.scala 206:34]
  wire  cout_3254 = cout_3170 & cout_3171; // @[Mul.scala 207:34]
  wire  sum_3255 = sum_3174 ^ sum_3175; // @[Mul.scala 206:34]
  wire  cout_3255 = sum_3174 & sum_3175; // @[Mul.scala 207:34]
  wire  sum_3256 = cout_3172 ^ cout_3173; // @[Mul.scala 206:34]
  wire  cout_3256 = cout_3172 & cout_3173; // @[Mul.scala 207:34]
  wire  sum_3257 = sum_3176 ^ sum_3177; // @[Mul.scala 206:34]
  wire  cout_3257 = sum_3176 & sum_3177; // @[Mul.scala 207:34]
  wire  sum_3258 = cout_3174 ^ cout_3175; // @[Mul.scala 206:34]
  wire  cout_3258 = cout_3174 & cout_3175; // @[Mul.scala 207:34]
  wire  sum_3259 = sum_3178 ^ sum_3179; // @[Mul.scala 206:34]
  wire  cout_3259 = sum_3178 & sum_3179; // @[Mul.scala 207:34]
  wire  sum_3260 = cout_3176 ^ cout_3177; // @[Mul.scala 206:34]
  wire  cout_3260 = cout_3176 & cout_3177; // @[Mul.scala 207:34]
  wire  sum_3261 = sum_3180 ^ sum_3181; // @[Mul.scala 206:34]
  wire  cout_3261 = sum_3180 & sum_3181; // @[Mul.scala 207:34]
  wire  sum_3262 = cout_3178 ^ cout_3179; // @[Mul.scala 206:34]
  wire  cout_3262 = cout_3178 & cout_3179; // @[Mul.scala 207:34]
  wire  sum_3263 = sum_3182 ^ sum_3183; // @[Mul.scala 206:34]
  wire  cout_3263 = sum_3182 & sum_3183; // @[Mul.scala 207:34]
  wire  sum_3264 = cout_3180 ^ cout_3181; // @[Mul.scala 206:34]
  wire  cout_3264 = cout_3180 & cout_3181; // @[Mul.scala 207:34]
  wire  sum_3265 = sum_3184 ^ sum_3185; // @[Mul.scala 206:34]
  wire  cout_3265 = sum_3184 & sum_3185; // @[Mul.scala 207:34]
  wire  sum_3266 = cout_3182 ^ cout_3183; // @[Mul.scala 206:34]
  wire  cout_3266 = cout_3182 & cout_3183; // @[Mul.scala 207:34]
  wire  sum_3267 = sum_3186 ^ sum_3187; // @[Mul.scala 206:34]
  wire  cout_3267 = sum_3186 & sum_3187; // @[Mul.scala 207:34]
  wire  sum_3268 = cout_3184 ^ cout_3185; // @[Mul.scala 206:34]
  wire  cout_3268 = cout_3184 & cout_3185; // @[Mul.scala 207:34]
  wire  sum_3269 = sum_3188 ^ sum_3189; // @[Mul.scala 206:34]
  wire  cout_3269 = sum_3188 & sum_3189; // @[Mul.scala 207:34]
  wire  sum_3270 = cout_3186 ^ cout_3187; // @[Mul.scala 206:34]
  wire  cout_3270 = cout_3186 & cout_3187; // @[Mul.scala 207:34]
  wire  sum_3271 = sum_3190 ^ sum_3191; // @[Mul.scala 206:34]
  wire  cout_3271 = sum_3190 & sum_3191; // @[Mul.scala 207:34]
  wire  sum_3272 = cout_3188 ^ cout_3189; // @[Mul.scala 206:34]
  wire  cout_3272 = cout_3188 & cout_3189; // @[Mul.scala 207:34]
  wire  sum_3273 = sum_3192 ^ sum_3193; // @[Mul.scala 206:34]
  wire  cout_3273 = sum_3192 & sum_3193; // @[Mul.scala 207:34]
  wire  sum_3274 = cout_3190 ^ cout_3191; // @[Mul.scala 206:34]
  wire  cout_3274 = cout_3190 & cout_3191; // @[Mul.scala 207:34]
  wire  sum_3275 = sum_3194 ^ sum_3195; // @[Mul.scala 206:34]
  wire  cout_3275 = sum_3194 & sum_3195; // @[Mul.scala 207:34]
  wire  sum_3276 = cout_3192 ^ cout_3193; // @[Mul.scala 206:34]
  wire  cout_3276 = cout_3192 & cout_3193; // @[Mul.scala 207:34]
  wire  sum_3277 = sum_3196 ^ sum_3197; // @[Mul.scala 206:34]
  wire  cout_3277 = sum_3196 & sum_3197; // @[Mul.scala 207:34]
  wire  sum_3278 = cout_3194 ^ cout_3195; // @[Mul.scala 206:34]
  wire  cout_3278 = cout_3194 & cout_3195; // @[Mul.scala 207:34]
  wire  sum_3279 = sum_3198 ^ sum_3199; // @[Mul.scala 206:34]
  wire  cout_3279 = sum_3198 & sum_3199; // @[Mul.scala 207:34]
  wire  sum_3280 = cout_3196 ^ cout_3197; // @[Mul.scala 206:34]
  wire  cout_3280 = cout_3196 & cout_3197; // @[Mul.scala 207:34]
  wire  sum_3281 = sum_3200 ^ sum_3201; // @[Mul.scala 206:34]
  wire  cout_3281 = sum_3200 & sum_3201; // @[Mul.scala 207:34]
  wire  sum_3282 = cout_3198 ^ cout_3199; // @[Mul.scala 206:34]
  wire  cout_3282 = cout_3198 & cout_3199; // @[Mul.scala 207:34]
  wire  sum_3283 = sum_3202 ^ sum_3203; // @[Mul.scala 206:34]
  wire  cout_3283 = sum_3202 & sum_3203; // @[Mul.scala 207:34]
  wire  sum_3284 = cout_3200 ^ cout_3201; // @[Mul.scala 206:34]
  wire  cout_3284 = cout_3200 & cout_3201; // @[Mul.scala 207:34]
  wire  _sum_T_3953 = sum_3204 ^ cout_3202; // @[Mul.scala 191:34]
  wire  sum_3285 = sum_3204 ^ cout_3202 ^ cout_3203; // @[Mul.scala 191:42]
  wire  cout_3285 = sum_3204 & cout_3202 | _sum_T_3953 & cout_3203; // @[Mul.scala 192:44]
  wire  sum_3286 = sum_3205 ^ cout_3204; // @[Mul.scala 206:34]
  wire  cout_3286 = sum_3205 & cout_3204; // @[Mul.scala 207:34]
  wire  sum_3287 = sum_3206 ^ cout_3205; // @[Mul.scala 206:34]
  wire  cout_3287 = sum_3206 & cout_3205; // @[Mul.scala 207:34]
  wire  sum_3288 = sum_3207 ^ cout_3206; // @[Mul.scala 206:34]
  wire  cout_3288 = sum_3207 & cout_3206; // @[Mul.scala 207:34]
  wire  sum_3289 = sum_3208 ^ cout_3207; // @[Mul.scala 206:34]
  wire  cout_3289 = sum_3208 & cout_3207; // @[Mul.scala 207:34]
  wire  sum_3290 = sum_3209 ^ cout_3208; // @[Mul.scala 206:34]
  wire  sum_3327 = sum_3246 ^ cout_3245; // @[Mul.scala 206:34]
  wire  cout_3327 = sum_3246 & cout_3245; // @[Mul.scala 207:34]
  wire  sum_3328 = sum_3247 ^ cout_3246; // @[Mul.scala 206:34]
  wire  cout_3328 = sum_3247 & cout_3246; // @[Mul.scala 207:34]
  wire  sum_3329 = sum_3248 ^ cout_3247; // @[Mul.scala 206:34]
  wire  cout_3329 = sum_3248 & cout_3247; // @[Mul.scala 207:34]
  wire  _sum_T_3999 = sum_3249 ^ sum_3250; // @[Mul.scala 191:34]
  wire  sum_3330 = sum_3249 ^ sum_3250 ^ cout_3248; // @[Mul.scala 191:42]
  wire  cout_3330 = sum_3249 & sum_3250 | _sum_T_3999 & cout_3248; // @[Mul.scala 192:44]
  wire  sum_3331 = sum_3251 ^ sum_3252; // @[Mul.scala 206:34]
  wire  cout_3331 = sum_3251 & sum_3252; // @[Mul.scala 207:34]
  wire  sum_3332 = cout_3249 ^ cout_3250; // @[Mul.scala 206:34]
  wire  cout_3332 = cout_3249 & cout_3250; // @[Mul.scala 207:34]
  wire  sum_3333 = sum_3253 ^ sum_3254; // @[Mul.scala 206:34]
  wire  cout_3333 = sum_3253 & sum_3254; // @[Mul.scala 207:34]
  wire  sum_3334 = cout_3251 ^ cout_3252; // @[Mul.scala 206:34]
  wire  cout_3334 = cout_3251 & cout_3252; // @[Mul.scala 207:34]
  wire  sum_3335 = sum_3255 ^ sum_3256; // @[Mul.scala 206:34]
  wire  cout_3335 = sum_3255 & sum_3256; // @[Mul.scala 207:34]
  wire  sum_3336 = cout_3253 ^ cout_3254; // @[Mul.scala 206:34]
  wire  cout_3336 = cout_3253 & cout_3254; // @[Mul.scala 207:34]
  wire  sum_3337 = sum_3257 ^ sum_3258; // @[Mul.scala 206:34]
  wire  cout_3337 = sum_3257 & sum_3258; // @[Mul.scala 207:34]
  wire  sum_3338 = cout_3255 ^ cout_3256; // @[Mul.scala 206:34]
  wire  cout_3338 = cout_3255 & cout_3256; // @[Mul.scala 207:34]
  wire  sum_3339 = sum_3259 ^ sum_3260; // @[Mul.scala 206:34]
  wire  cout_3339 = sum_3259 & sum_3260; // @[Mul.scala 207:34]
  wire  sum_3340 = cout_3257 ^ cout_3258; // @[Mul.scala 206:34]
  wire  cout_3340 = cout_3257 & cout_3258; // @[Mul.scala 207:34]
  wire  sum_3341 = sum_3261 ^ sum_3262; // @[Mul.scala 206:34]
  wire  cout_3341 = sum_3261 & sum_3262; // @[Mul.scala 207:34]
  wire  sum_3342 = cout_3259 ^ cout_3260; // @[Mul.scala 206:34]
  wire  cout_3342 = cout_3259 & cout_3260; // @[Mul.scala 207:34]
  wire  sum_3343 = sum_3263 ^ sum_3264; // @[Mul.scala 206:34]
  wire  cout_3343 = sum_3263 & sum_3264; // @[Mul.scala 207:34]
  wire  sum_3344 = cout_3261 ^ cout_3262; // @[Mul.scala 206:34]
  wire  cout_3344 = cout_3261 & cout_3262; // @[Mul.scala 207:34]
  wire  sum_3345 = sum_3265 ^ sum_3266; // @[Mul.scala 206:34]
  wire  cout_3345 = sum_3265 & sum_3266; // @[Mul.scala 207:34]
  wire  sum_3346 = cout_3263 ^ cout_3264; // @[Mul.scala 206:34]
  wire  cout_3346 = cout_3263 & cout_3264; // @[Mul.scala 207:34]
  wire  sum_3347 = sum_3267 ^ sum_3268; // @[Mul.scala 206:34]
  wire  cout_3347 = sum_3267 & sum_3268; // @[Mul.scala 207:34]
  wire  sum_3348 = cout_3265 ^ cout_3266; // @[Mul.scala 206:34]
  wire  cout_3348 = cout_3265 & cout_3266; // @[Mul.scala 207:34]
  wire  sum_3349 = sum_3269 ^ sum_3270; // @[Mul.scala 206:34]
  wire  cout_3349 = sum_3269 & sum_3270; // @[Mul.scala 207:34]
  wire  sum_3350 = cout_3267 ^ cout_3268; // @[Mul.scala 206:34]
  wire  cout_3350 = cout_3267 & cout_3268; // @[Mul.scala 207:34]
  wire  sum_3351 = sum_3271 ^ sum_3272; // @[Mul.scala 206:34]
  wire  cout_3351 = sum_3271 & sum_3272; // @[Mul.scala 207:34]
  wire  sum_3352 = cout_3269 ^ cout_3270; // @[Mul.scala 206:34]
  wire  cout_3352 = cout_3269 & cout_3270; // @[Mul.scala 207:34]
  wire  sum_3353 = sum_3273 ^ sum_3274; // @[Mul.scala 206:34]
  wire  cout_3353 = sum_3273 & sum_3274; // @[Mul.scala 207:34]
  wire  sum_3354 = cout_3271 ^ cout_3272; // @[Mul.scala 206:34]
  wire  cout_3354 = cout_3271 & cout_3272; // @[Mul.scala 207:34]
  wire  sum_3355 = sum_3275 ^ sum_3276; // @[Mul.scala 206:34]
  wire  cout_3355 = sum_3275 & sum_3276; // @[Mul.scala 207:34]
  wire  sum_3356 = cout_3273 ^ cout_3274; // @[Mul.scala 206:34]
  wire  cout_3356 = cout_3273 & cout_3274; // @[Mul.scala 207:34]
  wire  sum_3357 = sum_3277 ^ sum_3278; // @[Mul.scala 206:34]
  wire  cout_3357 = sum_3277 & sum_3278; // @[Mul.scala 207:34]
  wire  sum_3358 = cout_3275 ^ cout_3276; // @[Mul.scala 206:34]
  wire  cout_3358 = cout_3275 & cout_3276; // @[Mul.scala 207:34]
  wire  sum_3359 = sum_3279 ^ sum_3280; // @[Mul.scala 206:34]
  wire  cout_3359 = sum_3279 & sum_3280; // @[Mul.scala 207:34]
  wire  sum_3360 = cout_3277 ^ cout_3278; // @[Mul.scala 206:34]
  wire  cout_3360 = cout_3277 & cout_3278; // @[Mul.scala 207:34]
  wire  sum_3361 = sum_3281 ^ sum_3282; // @[Mul.scala 206:34]
  wire  cout_3361 = sum_3281 & sum_3282; // @[Mul.scala 207:34]
  wire  sum_3362 = cout_3279 ^ cout_3280; // @[Mul.scala 206:34]
  wire  cout_3362 = cout_3279 & cout_3280; // @[Mul.scala 207:34]
  wire  sum_3363 = sum_3283 ^ sum_3284; // @[Mul.scala 206:34]
  wire  cout_3363 = sum_3283 & sum_3284; // @[Mul.scala 207:34]
  wire  sum_3364 = cout_3281 ^ cout_3282; // @[Mul.scala 206:34]
  wire  cout_3364 = cout_3281 & cout_3282; // @[Mul.scala 207:34]
  wire  _sum_T_4035 = sum_3285 ^ cout_3283; // @[Mul.scala 191:34]
  wire  sum_3365 = sum_3285 ^ cout_3283 ^ cout_3284; // @[Mul.scala 191:42]
  wire  cout_3365 = sum_3285 & cout_3283 | _sum_T_4035 & cout_3284; // @[Mul.scala 192:44]
  wire  sum_3366 = sum_3286 ^ cout_3285; // @[Mul.scala 206:34]
  wire  cout_3366 = sum_3286 & cout_3285; // @[Mul.scala 207:34]
  wire  sum_3367 = sum_3287 ^ cout_3286; // @[Mul.scala 206:34]
  wire  cout_3367 = sum_3287 & cout_3286; // @[Mul.scala 207:34]
  wire  sum_3368 = sum_3288 ^ cout_3287; // @[Mul.scala 206:34]
  wire  cout_3368 = sum_3288 & cout_3287; // @[Mul.scala 207:34]
  wire  sum_3369 = sum_3289 ^ cout_3288; // @[Mul.scala 206:34]
  wire  cout_3369 = sum_3289 & cout_3288; // @[Mul.scala 207:34]
  wire  sum_3370 = sum_3290 ^ cout_3289; // @[Mul.scala 206:34]
  wire  sum_3408 = sum_3328 ^ cout_3327; // @[Mul.scala 206:34]
  wire  cout_3408 = sum_3328 & cout_3327; // @[Mul.scala 207:34]
  wire  sum_3409 = sum_3329 ^ cout_3328; // @[Mul.scala 206:34]
  wire  cout_3409 = sum_3329 & cout_3328; // @[Mul.scala 207:34]
  wire  sum_3410 = sum_3330 ^ cout_3329; // @[Mul.scala 206:34]
  wire  cout_3410 = sum_3330 & cout_3329; // @[Mul.scala 207:34]
  wire  _sum_T_4082 = sum_3331 ^ sum_3332; // @[Mul.scala 191:34]
  wire  sum_3411 = sum_3331 ^ sum_3332 ^ cout_3330; // @[Mul.scala 191:42]
  wire  cout_3411 = sum_3331 & sum_3332 | _sum_T_4082 & cout_3330; // @[Mul.scala 192:44]
  wire  sum_3412 = sum_3333 ^ sum_3334; // @[Mul.scala 206:34]
  wire  cout_3412 = sum_3333 & sum_3334; // @[Mul.scala 207:34]
  wire  sum_3413 = cout_3331 ^ cout_3332; // @[Mul.scala 206:34]
  wire  cout_3413 = cout_3331 & cout_3332; // @[Mul.scala 207:34]
  wire  sum_3414 = sum_3335 ^ sum_3336; // @[Mul.scala 206:34]
  wire  cout_3414 = sum_3335 & sum_3336; // @[Mul.scala 207:34]
  wire  sum_3415 = cout_3333 ^ cout_3334; // @[Mul.scala 206:34]
  wire  cout_3415 = cout_3333 & cout_3334; // @[Mul.scala 207:34]
  wire  sum_3416 = sum_3337 ^ sum_3338; // @[Mul.scala 206:34]
  wire  cout_3416 = sum_3337 & sum_3338; // @[Mul.scala 207:34]
  wire  sum_3417 = cout_3335 ^ cout_3336; // @[Mul.scala 206:34]
  wire  cout_3417 = cout_3335 & cout_3336; // @[Mul.scala 207:34]
  wire  sum_3418 = sum_3339 ^ sum_3340; // @[Mul.scala 206:34]
  wire  cout_3418 = sum_3339 & sum_3340; // @[Mul.scala 207:34]
  wire  sum_3419 = cout_3337 ^ cout_3338; // @[Mul.scala 206:34]
  wire  cout_3419 = cout_3337 & cout_3338; // @[Mul.scala 207:34]
  wire  sum_3420 = sum_3341 ^ sum_3342; // @[Mul.scala 206:34]
  wire  cout_3420 = sum_3341 & sum_3342; // @[Mul.scala 207:34]
  wire  sum_3421 = cout_3339 ^ cout_3340; // @[Mul.scala 206:34]
  wire  cout_3421 = cout_3339 & cout_3340; // @[Mul.scala 207:34]
  wire  sum_3422 = sum_3343 ^ sum_3344; // @[Mul.scala 206:34]
  wire  cout_3422 = sum_3343 & sum_3344; // @[Mul.scala 207:34]
  wire  sum_3423 = cout_3341 ^ cout_3342; // @[Mul.scala 206:34]
  wire  cout_3423 = cout_3341 & cout_3342; // @[Mul.scala 207:34]
  wire  sum_3424 = sum_3345 ^ sum_3346; // @[Mul.scala 206:34]
  wire  cout_3424 = sum_3345 & sum_3346; // @[Mul.scala 207:34]
  wire  sum_3425 = cout_3343 ^ cout_3344; // @[Mul.scala 206:34]
  wire  cout_3425 = cout_3343 & cout_3344; // @[Mul.scala 207:34]
  wire  sum_3426 = sum_3347 ^ sum_3348; // @[Mul.scala 206:34]
  wire  cout_3426 = sum_3347 & sum_3348; // @[Mul.scala 207:34]
  wire  sum_3427 = cout_3345 ^ cout_3346; // @[Mul.scala 206:34]
  wire  cout_3427 = cout_3345 & cout_3346; // @[Mul.scala 207:34]
  wire  sum_3428 = sum_3349 ^ sum_3350; // @[Mul.scala 206:34]
  wire  cout_3428 = sum_3349 & sum_3350; // @[Mul.scala 207:34]
  wire  sum_3429 = cout_3347 ^ cout_3348; // @[Mul.scala 206:34]
  wire  cout_3429 = cout_3347 & cout_3348; // @[Mul.scala 207:34]
  wire  sum_3430 = sum_3351 ^ sum_3352; // @[Mul.scala 206:34]
  wire  cout_3430 = sum_3351 & sum_3352; // @[Mul.scala 207:34]
  wire  sum_3431 = cout_3349 ^ cout_3350; // @[Mul.scala 206:34]
  wire  cout_3431 = cout_3349 & cout_3350; // @[Mul.scala 207:34]
  wire  sum_3432 = sum_3353 ^ sum_3354; // @[Mul.scala 206:34]
  wire  cout_3432 = sum_3353 & sum_3354; // @[Mul.scala 207:34]
  wire  sum_3433 = cout_3351 ^ cout_3352; // @[Mul.scala 206:34]
  wire  cout_3433 = cout_3351 & cout_3352; // @[Mul.scala 207:34]
  wire  sum_3434 = sum_3355 ^ sum_3356; // @[Mul.scala 206:34]
  wire  cout_3434 = sum_3355 & sum_3356; // @[Mul.scala 207:34]
  wire  sum_3435 = cout_3353 ^ cout_3354; // @[Mul.scala 206:34]
  wire  cout_3435 = cout_3353 & cout_3354; // @[Mul.scala 207:34]
  wire  sum_3436 = sum_3357 ^ sum_3358; // @[Mul.scala 206:34]
  wire  cout_3436 = sum_3357 & sum_3358; // @[Mul.scala 207:34]
  wire  sum_3437 = cout_3355 ^ cout_3356; // @[Mul.scala 206:34]
  wire  cout_3437 = cout_3355 & cout_3356; // @[Mul.scala 207:34]
  wire  sum_3438 = sum_3359 ^ sum_3360; // @[Mul.scala 206:34]
  wire  cout_3438 = sum_3359 & sum_3360; // @[Mul.scala 207:34]
  wire  sum_3439 = cout_3357 ^ cout_3358; // @[Mul.scala 206:34]
  wire  cout_3439 = cout_3357 & cout_3358; // @[Mul.scala 207:34]
  wire  sum_3440 = sum_3361 ^ sum_3362; // @[Mul.scala 206:34]
  wire  cout_3440 = sum_3361 & sum_3362; // @[Mul.scala 207:34]
  wire  sum_3441 = cout_3359 ^ cout_3360; // @[Mul.scala 206:34]
  wire  cout_3441 = cout_3359 & cout_3360; // @[Mul.scala 207:34]
  wire  sum_3442 = sum_3363 ^ sum_3364; // @[Mul.scala 206:34]
  wire  cout_3442 = sum_3363 & sum_3364; // @[Mul.scala 207:34]
  wire  sum_3443 = cout_3361 ^ cout_3362; // @[Mul.scala 206:34]
  wire  cout_3443 = cout_3361 & cout_3362; // @[Mul.scala 207:34]
  wire  _sum_T_4116 = sum_3365 ^ cout_3363; // @[Mul.scala 191:34]
  wire  sum_3444 = sum_3365 ^ cout_3363 ^ cout_3364; // @[Mul.scala 191:42]
  wire  cout_3444 = sum_3365 & cout_3363 | _sum_T_4116 & cout_3364; // @[Mul.scala 192:44]
  wire  sum_3445 = sum_3366 ^ cout_3365; // @[Mul.scala 206:34]
  wire  cout_3445 = sum_3366 & cout_3365; // @[Mul.scala 207:34]
  wire  sum_3446 = sum_3367 ^ cout_3366; // @[Mul.scala 206:34]
  wire  cout_3446 = sum_3367 & cout_3366; // @[Mul.scala 207:34]
  wire  sum_3447 = sum_3368 ^ cout_3367; // @[Mul.scala 206:34]
  wire  cout_3447 = sum_3368 & cout_3367; // @[Mul.scala 207:34]
  wire  sum_3448 = sum_3369 ^ cout_3368; // @[Mul.scala 206:34]
  wire  cout_3448 = sum_3369 & cout_3368; // @[Mul.scala 207:34]
  wire  sum_3449 = sum_3370 ^ cout_3369; // @[Mul.scala 206:34]
  wire  sum_3488 = sum_3409 ^ cout_3408; // @[Mul.scala 206:34]
  wire  cout_3488 = sum_3409 & cout_3408; // @[Mul.scala 207:34]
  wire  sum_3489 = sum_3410 ^ cout_3409; // @[Mul.scala 206:34]
  wire  cout_3489 = sum_3410 & cout_3409; // @[Mul.scala 207:34]
  wire  sum_3490 = sum_3411 ^ cout_3410; // @[Mul.scala 206:34]
  wire  cout_3490 = sum_3411 & cout_3410; // @[Mul.scala 207:34]
  wire  _sum_T_4164 = sum_3412 ^ sum_3413; // @[Mul.scala 191:34]
  wire  sum_3491 = sum_3412 ^ sum_3413 ^ cout_3411; // @[Mul.scala 191:42]
  wire  cout_3491 = sum_3412 & sum_3413 | _sum_T_4164 & cout_3411; // @[Mul.scala 192:44]
  wire  sum_3492 = sum_3414 ^ sum_3415; // @[Mul.scala 206:34]
  wire  cout_3492 = sum_3414 & sum_3415; // @[Mul.scala 207:34]
  wire  sum_3493 = cout_3412 ^ cout_3413; // @[Mul.scala 206:34]
  wire  cout_3493 = cout_3412 & cout_3413; // @[Mul.scala 207:34]
  wire  sum_3494 = sum_3416 ^ sum_3417; // @[Mul.scala 206:34]
  wire  cout_3494 = sum_3416 & sum_3417; // @[Mul.scala 207:34]
  wire  sum_3495 = cout_3414 ^ cout_3415; // @[Mul.scala 206:34]
  wire  cout_3495 = cout_3414 & cout_3415; // @[Mul.scala 207:34]
  wire  sum_3496 = sum_3418 ^ sum_3419; // @[Mul.scala 206:34]
  wire  cout_3496 = sum_3418 & sum_3419; // @[Mul.scala 207:34]
  wire  sum_3497 = cout_3416 ^ cout_3417; // @[Mul.scala 206:34]
  wire  cout_3497 = cout_3416 & cout_3417; // @[Mul.scala 207:34]
  wire  sum_3498 = sum_3420 ^ sum_3421; // @[Mul.scala 206:34]
  wire  cout_3498 = sum_3420 & sum_3421; // @[Mul.scala 207:34]
  wire  sum_3499 = cout_3418 ^ cout_3419; // @[Mul.scala 206:34]
  wire  cout_3499 = cout_3418 & cout_3419; // @[Mul.scala 207:34]
  wire  sum_3500 = sum_3422 ^ sum_3423; // @[Mul.scala 206:34]
  wire  cout_3500 = sum_3422 & sum_3423; // @[Mul.scala 207:34]
  wire  sum_3501 = cout_3420 ^ cout_3421; // @[Mul.scala 206:34]
  wire  cout_3501 = cout_3420 & cout_3421; // @[Mul.scala 207:34]
  wire  sum_3502 = sum_3424 ^ sum_3425; // @[Mul.scala 206:34]
  wire  cout_3502 = sum_3424 & sum_3425; // @[Mul.scala 207:34]
  wire  sum_3503 = cout_3422 ^ cout_3423; // @[Mul.scala 206:34]
  wire  cout_3503 = cout_3422 & cout_3423; // @[Mul.scala 207:34]
  wire  sum_3504 = sum_3426 ^ sum_3427; // @[Mul.scala 206:34]
  wire  cout_3504 = sum_3426 & sum_3427; // @[Mul.scala 207:34]
  wire  sum_3505 = cout_3424 ^ cout_3425; // @[Mul.scala 206:34]
  wire  cout_3505 = cout_3424 & cout_3425; // @[Mul.scala 207:34]
  wire  sum_3506 = sum_3428 ^ sum_3429; // @[Mul.scala 206:34]
  wire  cout_3506 = sum_3428 & sum_3429; // @[Mul.scala 207:34]
  wire  sum_3507 = cout_3426 ^ cout_3427; // @[Mul.scala 206:34]
  wire  cout_3507 = cout_3426 & cout_3427; // @[Mul.scala 207:34]
  wire  sum_3508 = sum_3430 ^ sum_3431; // @[Mul.scala 206:34]
  wire  cout_3508 = sum_3430 & sum_3431; // @[Mul.scala 207:34]
  wire  sum_3509 = cout_3428 ^ cout_3429; // @[Mul.scala 206:34]
  wire  cout_3509 = cout_3428 & cout_3429; // @[Mul.scala 207:34]
  wire  sum_3510 = sum_3432 ^ sum_3433; // @[Mul.scala 206:34]
  wire  cout_3510 = sum_3432 & sum_3433; // @[Mul.scala 207:34]
  wire  sum_3511 = cout_3430 ^ cout_3431; // @[Mul.scala 206:34]
  wire  cout_3511 = cout_3430 & cout_3431; // @[Mul.scala 207:34]
  wire  sum_3512 = sum_3434 ^ sum_3435; // @[Mul.scala 206:34]
  wire  cout_3512 = sum_3434 & sum_3435; // @[Mul.scala 207:34]
  wire  sum_3513 = cout_3432 ^ cout_3433; // @[Mul.scala 206:34]
  wire  cout_3513 = cout_3432 & cout_3433; // @[Mul.scala 207:34]
  wire  sum_3514 = sum_3436 ^ sum_3437; // @[Mul.scala 206:34]
  wire  cout_3514 = sum_3436 & sum_3437; // @[Mul.scala 207:34]
  wire  sum_3515 = cout_3434 ^ cout_3435; // @[Mul.scala 206:34]
  wire  cout_3515 = cout_3434 & cout_3435; // @[Mul.scala 207:34]
  wire  sum_3516 = sum_3438 ^ sum_3439; // @[Mul.scala 206:34]
  wire  cout_3516 = sum_3438 & sum_3439; // @[Mul.scala 207:34]
  wire  sum_3517 = cout_3436 ^ cout_3437; // @[Mul.scala 206:34]
  wire  cout_3517 = cout_3436 & cout_3437; // @[Mul.scala 207:34]
  wire  sum_3518 = sum_3440 ^ sum_3441; // @[Mul.scala 206:34]
  wire  cout_3518 = sum_3440 & sum_3441; // @[Mul.scala 207:34]
  wire  sum_3519 = cout_3438 ^ cout_3439; // @[Mul.scala 206:34]
  wire  cout_3519 = cout_3438 & cout_3439; // @[Mul.scala 207:34]
  wire  sum_3520 = sum_3442 ^ sum_3443; // @[Mul.scala 206:34]
  wire  cout_3520 = sum_3442 & sum_3443; // @[Mul.scala 207:34]
  wire  sum_3521 = cout_3440 ^ cout_3441; // @[Mul.scala 206:34]
  wire  cout_3521 = cout_3440 & cout_3441; // @[Mul.scala 207:34]
  wire  _sum_T_4196 = sum_3444 ^ cout_3442; // @[Mul.scala 191:34]
  wire  sum_3522 = sum_3444 ^ cout_3442 ^ cout_3443; // @[Mul.scala 191:42]
  wire  cout_3522 = sum_3444 & cout_3442 | _sum_T_4196 & cout_3443; // @[Mul.scala 192:44]
  wire  sum_3523 = sum_3445 ^ cout_3444; // @[Mul.scala 206:34]
  wire  cout_3523 = sum_3445 & cout_3444; // @[Mul.scala 207:34]
  wire  sum_3524 = sum_3446 ^ cout_3445; // @[Mul.scala 206:34]
  wire  cout_3524 = sum_3446 & cout_3445; // @[Mul.scala 207:34]
  wire  sum_3525 = sum_3447 ^ cout_3446; // @[Mul.scala 206:34]
  wire  cout_3525 = sum_3447 & cout_3446; // @[Mul.scala 207:34]
  wire  sum_3526 = sum_3448 ^ cout_3447; // @[Mul.scala 206:34]
  wire  cout_3526 = sum_3448 & cout_3447; // @[Mul.scala 207:34]
  wire  sum_3527 = sum_3449 ^ cout_3448; // @[Mul.scala 206:34]
  wire  sum_3567 = sum_3489 ^ cout_3488; // @[Mul.scala 206:34]
  wire  cout_3567 = sum_3489 & cout_3488; // @[Mul.scala 207:34]
  wire  sum_3568 = sum_3490 ^ cout_3489; // @[Mul.scala 206:34]
  wire  cout_3568 = sum_3490 & cout_3489; // @[Mul.scala 207:34]
  wire  sum_3569 = sum_3491 ^ cout_3490; // @[Mul.scala 206:34]
  wire  cout_3569 = sum_3491 & cout_3490; // @[Mul.scala 207:34]
  wire  _sum_T_4245 = sum_3492 ^ sum_3493; // @[Mul.scala 191:34]
  wire  sum_3570 = sum_3492 ^ sum_3493 ^ cout_3491; // @[Mul.scala 191:42]
  wire  cout_3570 = sum_3492 & sum_3493 | _sum_T_4245 & cout_3491; // @[Mul.scala 192:44]
  wire  sum_3571 = sum_3494 ^ sum_3495; // @[Mul.scala 206:34]
  wire  cout_3571 = sum_3494 & sum_3495; // @[Mul.scala 207:34]
  wire  sum_3572 = cout_3492 ^ cout_3493; // @[Mul.scala 206:34]
  wire  cout_3572 = cout_3492 & cout_3493; // @[Mul.scala 207:34]
  wire  sum_3573 = sum_3496 ^ sum_3497; // @[Mul.scala 206:34]
  wire  cout_3573 = sum_3496 & sum_3497; // @[Mul.scala 207:34]
  wire  sum_3574 = cout_3494 ^ cout_3495; // @[Mul.scala 206:34]
  wire  cout_3574 = cout_3494 & cout_3495; // @[Mul.scala 207:34]
  wire  sum_3575 = sum_3498 ^ sum_3499; // @[Mul.scala 206:34]
  wire  cout_3575 = sum_3498 & sum_3499; // @[Mul.scala 207:34]
  wire  sum_3576 = cout_3496 ^ cout_3497; // @[Mul.scala 206:34]
  wire  cout_3576 = cout_3496 & cout_3497; // @[Mul.scala 207:34]
  wire  sum_3577 = sum_3500 ^ sum_3501; // @[Mul.scala 206:34]
  wire  cout_3577 = sum_3500 & sum_3501; // @[Mul.scala 207:34]
  wire  sum_3578 = cout_3498 ^ cout_3499; // @[Mul.scala 206:34]
  wire  cout_3578 = cout_3498 & cout_3499; // @[Mul.scala 207:34]
  wire  sum_3579 = sum_3502 ^ sum_3503; // @[Mul.scala 206:34]
  wire  cout_3579 = sum_3502 & sum_3503; // @[Mul.scala 207:34]
  wire  sum_3580 = cout_3500 ^ cout_3501; // @[Mul.scala 206:34]
  wire  cout_3580 = cout_3500 & cout_3501; // @[Mul.scala 207:34]
  wire  sum_3581 = sum_3504 ^ sum_3505; // @[Mul.scala 206:34]
  wire  cout_3581 = sum_3504 & sum_3505; // @[Mul.scala 207:34]
  wire  sum_3582 = cout_3502 ^ cout_3503; // @[Mul.scala 206:34]
  wire  cout_3582 = cout_3502 & cout_3503; // @[Mul.scala 207:34]
  wire  sum_3583 = sum_3506 ^ sum_3507; // @[Mul.scala 206:34]
  wire  cout_3583 = sum_3506 & sum_3507; // @[Mul.scala 207:34]
  wire  sum_3584 = cout_3504 ^ cout_3505; // @[Mul.scala 206:34]
  wire  cout_3584 = cout_3504 & cout_3505; // @[Mul.scala 207:34]
  wire  sum_3585 = sum_3508 ^ sum_3509; // @[Mul.scala 206:34]
  wire  cout_3585 = sum_3508 & sum_3509; // @[Mul.scala 207:34]
  wire  sum_3586 = cout_3506 ^ cout_3507; // @[Mul.scala 206:34]
  wire  cout_3586 = cout_3506 & cout_3507; // @[Mul.scala 207:34]
  wire  sum_3587 = sum_3510 ^ sum_3511; // @[Mul.scala 206:34]
  wire  cout_3587 = sum_3510 & sum_3511; // @[Mul.scala 207:34]
  wire  sum_3588 = cout_3508 ^ cout_3509; // @[Mul.scala 206:34]
  wire  cout_3588 = cout_3508 & cout_3509; // @[Mul.scala 207:34]
  wire  sum_3589 = sum_3512 ^ sum_3513; // @[Mul.scala 206:34]
  wire  cout_3589 = sum_3512 & sum_3513; // @[Mul.scala 207:34]
  wire  sum_3590 = cout_3510 ^ cout_3511; // @[Mul.scala 206:34]
  wire  cout_3590 = cout_3510 & cout_3511; // @[Mul.scala 207:34]
  wire  sum_3591 = sum_3514 ^ sum_3515; // @[Mul.scala 206:34]
  wire  cout_3591 = sum_3514 & sum_3515; // @[Mul.scala 207:34]
  wire  sum_3592 = cout_3512 ^ cout_3513; // @[Mul.scala 206:34]
  wire  cout_3592 = cout_3512 & cout_3513; // @[Mul.scala 207:34]
  wire  sum_3593 = sum_3516 ^ sum_3517; // @[Mul.scala 206:34]
  wire  cout_3593 = sum_3516 & sum_3517; // @[Mul.scala 207:34]
  wire  sum_3594 = cout_3514 ^ cout_3515; // @[Mul.scala 206:34]
  wire  cout_3594 = cout_3514 & cout_3515; // @[Mul.scala 207:34]
  wire  sum_3595 = sum_3518 ^ sum_3519; // @[Mul.scala 206:34]
  wire  cout_3595 = sum_3518 & sum_3519; // @[Mul.scala 207:34]
  wire  sum_3596 = cout_3516 ^ cout_3517; // @[Mul.scala 206:34]
  wire  cout_3596 = cout_3516 & cout_3517; // @[Mul.scala 207:34]
  wire  sum_3597 = sum_3520 ^ sum_3521; // @[Mul.scala 206:34]
  wire  cout_3597 = sum_3520 & sum_3521; // @[Mul.scala 207:34]
  wire  sum_3598 = cout_3518 ^ cout_3519; // @[Mul.scala 206:34]
  wire  cout_3598 = cout_3518 & cout_3519; // @[Mul.scala 207:34]
  wire  _sum_T_4275 = sum_3522 ^ cout_3520; // @[Mul.scala 191:34]
  wire  sum_3599 = sum_3522 ^ cout_3520 ^ cout_3521; // @[Mul.scala 191:42]
  wire  cout_3599 = sum_3522 & cout_3520 | _sum_T_4275 & cout_3521; // @[Mul.scala 192:44]
  wire  sum_3600 = sum_3523 ^ cout_3522; // @[Mul.scala 206:34]
  wire  cout_3600 = sum_3523 & cout_3522; // @[Mul.scala 207:34]
  wire  sum_3601 = sum_3524 ^ cout_3523; // @[Mul.scala 206:34]
  wire  cout_3601 = sum_3524 & cout_3523; // @[Mul.scala 207:34]
  wire  sum_3602 = sum_3525 ^ cout_3524; // @[Mul.scala 206:34]
  wire  cout_3602 = sum_3525 & cout_3524; // @[Mul.scala 207:34]
  wire  sum_3603 = sum_3526 ^ cout_3525; // @[Mul.scala 206:34]
  wire  cout_3603 = sum_3526 & cout_3525; // @[Mul.scala 207:34]
  wire  sum_3604 = sum_3527 ^ cout_3526; // @[Mul.scala 206:34]
  wire  sum_3645 = sum_3568 ^ cout_3567; // @[Mul.scala 206:34]
  wire  cout_3645 = sum_3568 & cout_3567; // @[Mul.scala 207:34]
  wire  sum_3646 = sum_3569 ^ cout_3568; // @[Mul.scala 206:34]
  wire  cout_3646 = sum_3569 & cout_3568; // @[Mul.scala 207:34]
  wire  sum_3647 = sum_3570 ^ cout_3569; // @[Mul.scala 206:34]
  wire  cout_3647 = sum_3570 & cout_3569; // @[Mul.scala 207:34]
  wire  _sum_T_4325 = sum_3571 ^ sum_3572; // @[Mul.scala 191:34]
  wire  sum_3648 = sum_3571 ^ sum_3572 ^ cout_3570; // @[Mul.scala 191:42]
  wire  cout_3648 = sum_3571 & sum_3572 | _sum_T_4325 & cout_3570; // @[Mul.scala 192:44]
  wire  sum_3649 = sum_3573 ^ sum_3574; // @[Mul.scala 206:34]
  wire  cout_3649 = sum_3573 & sum_3574; // @[Mul.scala 207:34]
  wire  sum_3650 = cout_3571 ^ cout_3572; // @[Mul.scala 206:34]
  wire  cout_3650 = cout_3571 & cout_3572; // @[Mul.scala 207:34]
  wire  sum_3651 = sum_3575 ^ sum_3576; // @[Mul.scala 206:34]
  wire  cout_3651 = sum_3575 & sum_3576; // @[Mul.scala 207:34]
  wire  sum_3652 = cout_3573 ^ cout_3574; // @[Mul.scala 206:34]
  wire  cout_3652 = cout_3573 & cout_3574; // @[Mul.scala 207:34]
  wire  sum_3653 = sum_3577 ^ sum_3578; // @[Mul.scala 206:34]
  wire  cout_3653 = sum_3577 & sum_3578; // @[Mul.scala 207:34]
  wire  sum_3654 = cout_3575 ^ cout_3576; // @[Mul.scala 206:34]
  wire  cout_3654 = cout_3575 & cout_3576; // @[Mul.scala 207:34]
  wire  sum_3655 = sum_3579 ^ sum_3580; // @[Mul.scala 206:34]
  wire  cout_3655 = sum_3579 & sum_3580; // @[Mul.scala 207:34]
  wire  sum_3656 = cout_3577 ^ cout_3578; // @[Mul.scala 206:34]
  wire  cout_3656 = cout_3577 & cout_3578; // @[Mul.scala 207:34]
  wire  sum_3657 = sum_3581 ^ sum_3582; // @[Mul.scala 206:34]
  wire  cout_3657 = sum_3581 & sum_3582; // @[Mul.scala 207:34]
  wire  sum_3658 = cout_3579 ^ cout_3580; // @[Mul.scala 206:34]
  wire  cout_3658 = cout_3579 & cout_3580; // @[Mul.scala 207:34]
  wire  sum_3659 = sum_3583 ^ sum_3584; // @[Mul.scala 206:34]
  wire  cout_3659 = sum_3583 & sum_3584; // @[Mul.scala 207:34]
  wire  sum_3660 = cout_3581 ^ cout_3582; // @[Mul.scala 206:34]
  wire  cout_3660 = cout_3581 & cout_3582; // @[Mul.scala 207:34]
  wire  sum_3661 = sum_3585 ^ sum_3586; // @[Mul.scala 206:34]
  wire  cout_3661 = sum_3585 & sum_3586; // @[Mul.scala 207:34]
  wire  sum_3662 = cout_3583 ^ cout_3584; // @[Mul.scala 206:34]
  wire  cout_3662 = cout_3583 & cout_3584; // @[Mul.scala 207:34]
  wire  sum_3663 = sum_3587 ^ sum_3588; // @[Mul.scala 206:34]
  wire  cout_3663 = sum_3587 & sum_3588; // @[Mul.scala 207:34]
  wire  sum_3664 = cout_3585 ^ cout_3586; // @[Mul.scala 206:34]
  wire  cout_3664 = cout_3585 & cout_3586; // @[Mul.scala 207:34]
  wire  sum_3665 = sum_3589 ^ sum_3590; // @[Mul.scala 206:34]
  wire  cout_3665 = sum_3589 & sum_3590; // @[Mul.scala 207:34]
  wire  sum_3666 = cout_3587 ^ cout_3588; // @[Mul.scala 206:34]
  wire  cout_3666 = cout_3587 & cout_3588; // @[Mul.scala 207:34]
  wire  sum_3667 = sum_3591 ^ sum_3592; // @[Mul.scala 206:34]
  wire  cout_3667 = sum_3591 & sum_3592; // @[Mul.scala 207:34]
  wire  sum_3668 = cout_3589 ^ cout_3590; // @[Mul.scala 206:34]
  wire  cout_3668 = cout_3589 & cout_3590; // @[Mul.scala 207:34]
  wire  sum_3669 = sum_3593 ^ sum_3594; // @[Mul.scala 206:34]
  wire  cout_3669 = sum_3593 & sum_3594; // @[Mul.scala 207:34]
  wire  sum_3670 = cout_3591 ^ cout_3592; // @[Mul.scala 206:34]
  wire  cout_3670 = cout_3591 & cout_3592; // @[Mul.scala 207:34]
  wire  sum_3671 = sum_3595 ^ sum_3596; // @[Mul.scala 206:34]
  wire  cout_3671 = sum_3595 & sum_3596; // @[Mul.scala 207:34]
  wire  sum_3672 = cout_3593 ^ cout_3594; // @[Mul.scala 206:34]
  wire  cout_3672 = cout_3593 & cout_3594; // @[Mul.scala 207:34]
  wire  sum_3673 = sum_3597 ^ sum_3598; // @[Mul.scala 206:34]
  wire  cout_3673 = sum_3597 & sum_3598; // @[Mul.scala 207:34]
  wire  sum_3674 = cout_3595 ^ cout_3596; // @[Mul.scala 206:34]
  wire  cout_3674 = cout_3595 & cout_3596; // @[Mul.scala 207:34]
  wire  _sum_T_4353 = sum_3599 ^ cout_3597; // @[Mul.scala 191:34]
  wire  sum_3675 = sum_3599 ^ cout_3597 ^ cout_3598; // @[Mul.scala 191:42]
  wire  cout_3675 = sum_3599 & cout_3597 | _sum_T_4353 & cout_3598; // @[Mul.scala 192:44]
  wire  sum_3676 = sum_3600 ^ cout_3599; // @[Mul.scala 206:34]
  wire  cout_3676 = sum_3600 & cout_3599; // @[Mul.scala 207:34]
  wire  sum_3677 = sum_3601 ^ cout_3600; // @[Mul.scala 206:34]
  wire  cout_3677 = sum_3601 & cout_3600; // @[Mul.scala 207:34]
  wire  sum_3678 = sum_3602 ^ cout_3601; // @[Mul.scala 206:34]
  wire  cout_3678 = sum_3602 & cout_3601; // @[Mul.scala 207:34]
  wire  sum_3679 = sum_3603 ^ cout_3602; // @[Mul.scala 206:34]
  wire  cout_3679 = sum_3603 & cout_3602; // @[Mul.scala 207:34]
  wire  sum_3680 = sum_3604 ^ cout_3603; // @[Mul.scala 206:34]
  wire  sum_3722 = sum_3646 ^ cout_3645; // @[Mul.scala 206:34]
  wire  cout_3722 = sum_3646 & cout_3645; // @[Mul.scala 207:34]
  wire  sum_3723 = sum_3647 ^ cout_3646; // @[Mul.scala 206:34]
  wire  cout_3723 = sum_3647 & cout_3646; // @[Mul.scala 207:34]
  wire  sum_3724 = sum_3648 ^ cout_3647; // @[Mul.scala 206:34]
  wire  cout_3724 = sum_3648 & cout_3647; // @[Mul.scala 207:34]
  wire  _sum_T_4404 = sum_3649 ^ sum_3650; // @[Mul.scala 191:34]
  wire  sum_3725 = sum_3649 ^ sum_3650 ^ cout_3648; // @[Mul.scala 191:42]
  wire  cout_3725 = sum_3649 & sum_3650 | _sum_T_4404 & cout_3648; // @[Mul.scala 192:44]
  wire  sum_3726 = sum_3651 ^ sum_3652; // @[Mul.scala 206:34]
  wire  cout_3726 = sum_3651 & sum_3652; // @[Mul.scala 207:34]
  wire  sum_3727 = cout_3649 ^ cout_3650; // @[Mul.scala 206:34]
  wire  cout_3727 = cout_3649 & cout_3650; // @[Mul.scala 207:34]
  wire  sum_3728 = sum_3653 ^ sum_3654; // @[Mul.scala 206:34]
  wire  cout_3728 = sum_3653 & sum_3654; // @[Mul.scala 207:34]
  wire  sum_3729 = cout_3651 ^ cout_3652; // @[Mul.scala 206:34]
  wire  cout_3729 = cout_3651 & cout_3652; // @[Mul.scala 207:34]
  wire  sum_3730 = sum_3655 ^ sum_3656; // @[Mul.scala 206:34]
  wire  cout_3730 = sum_3655 & sum_3656; // @[Mul.scala 207:34]
  wire  sum_3731 = cout_3653 ^ cout_3654; // @[Mul.scala 206:34]
  wire  cout_3731 = cout_3653 & cout_3654; // @[Mul.scala 207:34]
  wire  sum_3732 = sum_3657 ^ sum_3658; // @[Mul.scala 206:34]
  wire  cout_3732 = sum_3657 & sum_3658; // @[Mul.scala 207:34]
  wire  sum_3733 = cout_3655 ^ cout_3656; // @[Mul.scala 206:34]
  wire  cout_3733 = cout_3655 & cout_3656; // @[Mul.scala 207:34]
  wire  sum_3734 = sum_3659 ^ sum_3660; // @[Mul.scala 206:34]
  wire  cout_3734 = sum_3659 & sum_3660; // @[Mul.scala 207:34]
  wire  sum_3735 = cout_3657 ^ cout_3658; // @[Mul.scala 206:34]
  wire  cout_3735 = cout_3657 & cout_3658; // @[Mul.scala 207:34]
  wire  sum_3736 = sum_3661 ^ sum_3662; // @[Mul.scala 206:34]
  wire  cout_3736 = sum_3661 & sum_3662; // @[Mul.scala 207:34]
  wire  sum_3737 = cout_3659 ^ cout_3660; // @[Mul.scala 206:34]
  wire  cout_3737 = cout_3659 & cout_3660; // @[Mul.scala 207:34]
  wire  sum_3738 = sum_3663 ^ sum_3664; // @[Mul.scala 206:34]
  wire  cout_3738 = sum_3663 & sum_3664; // @[Mul.scala 207:34]
  wire  sum_3739 = cout_3661 ^ cout_3662; // @[Mul.scala 206:34]
  wire  cout_3739 = cout_3661 & cout_3662; // @[Mul.scala 207:34]
  wire  sum_3740 = sum_3665 ^ sum_3666; // @[Mul.scala 206:34]
  wire  cout_3740 = sum_3665 & sum_3666; // @[Mul.scala 207:34]
  wire  sum_3741 = cout_3663 ^ cout_3664; // @[Mul.scala 206:34]
  wire  cout_3741 = cout_3663 & cout_3664; // @[Mul.scala 207:34]
  wire  sum_3742 = sum_3667 ^ sum_3668; // @[Mul.scala 206:34]
  wire  cout_3742 = sum_3667 & sum_3668; // @[Mul.scala 207:34]
  wire  sum_3743 = cout_3665 ^ cout_3666; // @[Mul.scala 206:34]
  wire  cout_3743 = cout_3665 & cout_3666; // @[Mul.scala 207:34]
  wire  sum_3744 = sum_3669 ^ sum_3670; // @[Mul.scala 206:34]
  wire  cout_3744 = sum_3669 & sum_3670; // @[Mul.scala 207:34]
  wire  sum_3745 = cout_3667 ^ cout_3668; // @[Mul.scala 206:34]
  wire  cout_3745 = cout_3667 & cout_3668; // @[Mul.scala 207:34]
  wire  sum_3746 = sum_3671 ^ sum_3672; // @[Mul.scala 206:34]
  wire  cout_3746 = sum_3671 & sum_3672; // @[Mul.scala 207:34]
  wire  sum_3747 = cout_3669 ^ cout_3670; // @[Mul.scala 206:34]
  wire  cout_3747 = cout_3669 & cout_3670; // @[Mul.scala 207:34]
  wire  sum_3748 = sum_3673 ^ sum_3674; // @[Mul.scala 206:34]
  wire  cout_3748 = sum_3673 & sum_3674; // @[Mul.scala 207:34]
  wire  sum_3749 = cout_3671 ^ cout_3672; // @[Mul.scala 206:34]
  wire  cout_3749 = cout_3671 & cout_3672; // @[Mul.scala 207:34]
  wire  _sum_T_4430 = sum_3675 ^ cout_3673; // @[Mul.scala 191:34]
  wire  sum_3750 = sum_3675 ^ cout_3673 ^ cout_3674; // @[Mul.scala 191:42]
  wire  cout_3750 = sum_3675 & cout_3673 | _sum_T_4430 & cout_3674; // @[Mul.scala 192:44]
  wire  sum_3751 = sum_3676 ^ cout_3675; // @[Mul.scala 206:34]
  wire  cout_3751 = sum_3676 & cout_3675; // @[Mul.scala 207:34]
  wire  sum_3752 = sum_3677 ^ cout_3676; // @[Mul.scala 206:34]
  wire  cout_3752 = sum_3677 & cout_3676; // @[Mul.scala 207:34]
  wire  sum_3753 = sum_3678 ^ cout_3677; // @[Mul.scala 206:34]
  wire  cout_3753 = sum_3678 & cout_3677; // @[Mul.scala 207:34]
  wire  sum_3754 = sum_3679 ^ cout_3678; // @[Mul.scala 206:34]
  wire  cout_3754 = sum_3679 & cout_3678; // @[Mul.scala 207:34]
  wire  sum_3755 = sum_3680 ^ cout_3679; // @[Mul.scala 206:34]
  wire  sum_3798 = sum_3723 ^ cout_3722; // @[Mul.scala 206:34]
  wire  cout_3798 = sum_3723 & cout_3722; // @[Mul.scala 207:34]
  wire  sum_3799 = sum_3724 ^ cout_3723; // @[Mul.scala 206:34]
  wire  cout_3799 = sum_3724 & cout_3723; // @[Mul.scala 207:34]
  wire  sum_3800 = sum_3725 ^ cout_3724; // @[Mul.scala 206:34]
  wire  cout_3800 = sum_3725 & cout_3724; // @[Mul.scala 207:34]
  wire  _sum_T_4482 = sum_3726 ^ sum_3727; // @[Mul.scala 191:34]
  wire  sum_3801 = sum_3726 ^ sum_3727 ^ cout_3725; // @[Mul.scala 191:42]
  wire  cout_3801 = sum_3726 & sum_3727 | _sum_T_4482 & cout_3725; // @[Mul.scala 192:44]
  wire  sum_3802 = sum_3728 ^ sum_3729; // @[Mul.scala 206:34]
  wire  cout_3802 = sum_3728 & sum_3729; // @[Mul.scala 207:34]
  wire  sum_3803 = cout_3726 ^ cout_3727; // @[Mul.scala 206:34]
  wire  cout_3803 = cout_3726 & cout_3727; // @[Mul.scala 207:34]
  wire  sum_3804 = sum_3730 ^ sum_3731; // @[Mul.scala 206:34]
  wire  cout_3804 = sum_3730 & sum_3731; // @[Mul.scala 207:34]
  wire  sum_3805 = cout_3728 ^ cout_3729; // @[Mul.scala 206:34]
  wire  cout_3805 = cout_3728 & cout_3729; // @[Mul.scala 207:34]
  wire  sum_3806 = sum_3732 ^ sum_3733; // @[Mul.scala 206:34]
  wire  cout_3806 = sum_3732 & sum_3733; // @[Mul.scala 207:34]
  wire  sum_3807 = cout_3730 ^ cout_3731; // @[Mul.scala 206:34]
  wire  cout_3807 = cout_3730 & cout_3731; // @[Mul.scala 207:34]
  wire  sum_3808 = sum_3734 ^ sum_3735; // @[Mul.scala 206:34]
  wire  cout_3808 = sum_3734 & sum_3735; // @[Mul.scala 207:34]
  wire  sum_3809 = cout_3732 ^ cout_3733; // @[Mul.scala 206:34]
  wire  cout_3809 = cout_3732 & cout_3733; // @[Mul.scala 207:34]
  wire  sum_3810 = sum_3736 ^ sum_3737; // @[Mul.scala 206:34]
  wire  cout_3810 = sum_3736 & sum_3737; // @[Mul.scala 207:34]
  wire  sum_3811 = cout_3734 ^ cout_3735; // @[Mul.scala 206:34]
  wire  cout_3811 = cout_3734 & cout_3735; // @[Mul.scala 207:34]
  wire  sum_3812 = sum_3738 ^ sum_3739; // @[Mul.scala 206:34]
  wire  cout_3812 = sum_3738 & sum_3739; // @[Mul.scala 207:34]
  wire  sum_3813 = cout_3736 ^ cout_3737; // @[Mul.scala 206:34]
  wire  cout_3813 = cout_3736 & cout_3737; // @[Mul.scala 207:34]
  wire  sum_3814 = sum_3740 ^ sum_3741; // @[Mul.scala 206:34]
  wire  cout_3814 = sum_3740 & sum_3741; // @[Mul.scala 207:34]
  wire  sum_3815 = cout_3738 ^ cout_3739; // @[Mul.scala 206:34]
  wire  cout_3815 = cout_3738 & cout_3739; // @[Mul.scala 207:34]
  wire  sum_3816 = sum_3742 ^ sum_3743; // @[Mul.scala 206:34]
  wire  cout_3816 = sum_3742 & sum_3743; // @[Mul.scala 207:34]
  wire  sum_3817 = cout_3740 ^ cout_3741; // @[Mul.scala 206:34]
  wire  cout_3817 = cout_3740 & cout_3741; // @[Mul.scala 207:34]
  wire  sum_3818 = sum_3744 ^ sum_3745; // @[Mul.scala 206:34]
  wire  cout_3818 = sum_3744 & sum_3745; // @[Mul.scala 207:34]
  wire  sum_3819 = cout_3742 ^ cout_3743; // @[Mul.scala 206:34]
  wire  cout_3819 = cout_3742 & cout_3743; // @[Mul.scala 207:34]
  wire  sum_3820 = sum_3746 ^ sum_3747; // @[Mul.scala 206:34]
  wire  cout_3820 = sum_3746 & sum_3747; // @[Mul.scala 207:34]
  wire  sum_3821 = cout_3744 ^ cout_3745; // @[Mul.scala 206:34]
  wire  cout_3821 = cout_3744 & cout_3745; // @[Mul.scala 207:34]
  wire  sum_3822 = sum_3748 ^ sum_3749; // @[Mul.scala 206:34]
  wire  cout_3822 = sum_3748 & sum_3749; // @[Mul.scala 207:34]
  wire  sum_3823 = cout_3746 ^ cout_3747; // @[Mul.scala 206:34]
  wire  cout_3823 = cout_3746 & cout_3747; // @[Mul.scala 207:34]
  wire  _sum_T_4506 = sum_3750 ^ cout_3748; // @[Mul.scala 191:34]
  wire  sum_3824 = sum_3750 ^ cout_3748 ^ cout_3749; // @[Mul.scala 191:42]
  wire  cout_3824 = sum_3750 & cout_3748 | _sum_T_4506 & cout_3749; // @[Mul.scala 192:44]
  wire  sum_3825 = sum_3751 ^ cout_3750; // @[Mul.scala 206:34]
  wire  cout_3825 = sum_3751 & cout_3750; // @[Mul.scala 207:34]
  wire  sum_3826 = sum_3752 ^ cout_3751; // @[Mul.scala 206:34]
  wire  cout_3826 = sum_3752 & cout_3751; // @[Mul.scala 207:34]
  wire  sum_3827 = sum_3753 ^ cout_3752; // @[Mul.scala 206:34]
  wire  cout_3827 = sum_3753 & cout_3752; // @[Mul.scala 207:34]
  wire  sum_3828 = sum_3754 ^ cout_3753; // @[Mul.scala 206:34]
  wire  cout_3828 = sum_3754 & cout_3753; // @[Mul.scala 207:34]
  wire  sum_3829 = sum_3755 ^ cout_3754; // @[Mul.scala 206:34]
  wire  sum_3873 = sum_3799 ^ cout_3798; // @[Mul.scala 206:34]
  wire  cout_3873 = sum_3799 & cout_3798; // @[Mul.scala 207:34]
  wire  sum_3874 = sum_3800 ^ cout_3799; // @[Mul.scala 206:34]
  wire  cout_3874 = sum_3800 & cout_3799; // @[Mul.scala 207:34]
  wire  sum_3875 = sum_3801 ^ cout_3800; // @[Mul.scala 206:34]
  wire  cout_3875 = sum_3801 & cout_3800; // @[Mul.scala 207:34]
  wire  _sum_T_4559 = sum_3802 ^ sum_3803; // @[Mul.scala 191:34]
  wire  sum_3876 = sum_3802 ^ sum_3803 ^ cout_3801; // @[Mul.scala 191:42]
  wire  cout_3876 = sum_3802 & sum_3803 | _sum_T_4559 & cout_3801; // @[Mul.scala 192:44]
  wire  sum_3877 = sum_3804 ^ sum_3805; // @[Mul.scala 206:34]
  wire  cout_3877 = sum_3804 & sum_3805; // @[Mul.scala 207:34]
  wire  sum_3878 = cout_3802 ^ cout_3803; // @[Mul.scala 206:34]
  wire  cout_3878 = cout_3802 & cout_3803; // @[Mul.scala 207:34]
  wire  sum_3879 = sum_3806 ^ sum_3807; // @[Mul.scala 206:34]
  wire  cout_3879 = sum_3806 & sum_3807; // @[Mul.scala 207:34]
  wire  sum_3880 = cout_3804 ^ cout_3805; // @[Mul.scala 206:34]
  wire  cout_3880 = cout_3804 & cout_3805; // @[Mul.scala 207:34]
  wire  sum_3881 = sum_3808 ^ sum_3809; // @[Mul.scala 206:34]
  wire  cout_3881 = sum_3808 & sum_3809; // @[Mul.scala 207:34]
  wire  sum_3882 = cout_3806 ^ cout_3807; // @[Mul.scala 206:34]
  wire  cout_3882 = cout_3806 & cout_3807; // @[Mul.scala 207:34]
  wire  sum_3883 = sum_3810 ^ sum_3811; // @[Mul.scala 206:34]
  wire  cout_3883 = sum_3810 & sum_3811; // @[Mul.scala 207:34]
  wire  sum_3884 = cout_3808 ^ cout_3809; // @[Mul.scala 206:34]
  wire  cout_3884 = cout_3808 & cout_3809; // @[Mul.scala 207:34]
  wire  sum_3885 = sum_3812 ^ sum_3813; // @[Mul.scala 206:34]
  wire  cout_3885 = sum_3812 & sum_3813; // @[Mul.scala 207:34]
  wire  sum_3886 = cout_3810 ^ cout_3811; // @[Mul.scala 206:34]
  wire  cout_3886 = cout_3810 & cout_3811; // @[Mul.scala 207:34]
  wire  sum_3887 = sum_3814 ^ sum_3815; // @[Mul.scala 206:34]
  wire  cout_3887 = sum_3814 & sum_3815; // @[Mul.scala 207:34]
  wire  sum_3888 = cout_3812 ^ cout_3813; // @[Mul.scala 206:34]
  wire  cout_3888 = cout_3812 & cout_3813; // @[Mul.scala 207:34]
  wire  sum_3889 = sum_3816 ^ sum_3817; // @[Mul.scala 206:34]
  wire  cout_3889 = sum_3816 & sum_3817; // @[Mul.scala 207:34]
  wire  sum_3890 = cout_3814 ^ cout_3815; // @[Mul.scala 206:34]
  wire  cout_3890 = cout_3814 & cout_3815; // @[Mul.scala 207:34]
  wire  sum_3891 = sum_3818 ^ sum_3819; // @[Mul.scala 206:34]
  wire  cout_3891 = sum_3818 & sum_3819; // @[Mul.scala 207:34]
  wire  sum_3892 = cout_3816 ^ cout_3817; // @[Mul.scala 206:34]
  wire  cout_3892 = cout_3816 & cout_3817; // @[Mul.scala 207:34]
  wire  sum_3893 = sum_3820 ^ sum_3821; // @[Mul.scala 206:34]
  wire  cout_3893 = sum_3820 & sum_3821; // @[Mul.scala 207:34]
  wire  sum_3894 = cout_3818 ^ cout_3819; // @[Mul.scala 206:34]
  wire  cout_3894 = cout_3818 & cout_3819; // @[Mul.scala 207:34]
  wire  sum_3895 = sum_3822 ^ sum_3823; // @[Mul.scala 206:34]
  wire  cout_3895 = sum_3822 & sum_3823; // @[Mul.scala 207:34]
  wire  sum_3896 = cout_3820 ^ cout_3821; // @[Mul.scala 206:34]
  wire  cout_3896 = cout_3820 & cout_3821; // @[Mul.scala 207:34]
  wire  _sum_T_4581 = sum_3824 ^ cout_3822; // @[Mul.scala 191:34]
  wire  sum_3897 = sum_3824 ^ cout_3822 ^ cout_3823; // @[Mul.scala 191:42]
  wire  cout_3897 = sum_3824 & cout_3822 | _sum_T_4581 & cout_3823; // @[Mul.scala 192:44]
  wire  sum_3898 = sum_3825 ^ cout_3824; // @[Mul.scala 206:34]
  wire  cout_3898 = sum_3825 & cout_3824; // @[Mul.scala 207:34]
  wire  sum_3899 = sum_3826 ^ cout_3825; // @[Mul.scala 206:34]
  wire  cout_3899 = sum_3826 & cout_3825; // @[Mul.scala 207:34]
  wire  sum_3900 = sum_3827 ^ cout_3826; // @[Mul.scala 206:34]
  wire  cout_3900 = sum_3827 & cout_3826; // @[Mul.scala 207:34]
  wire  sum_3901 = sum_3828 ^ cout_3827; // @[Mul.scala 206:34]
  wire  cout_3901 = sum_3828 & cout_3827; // @[Mul.scala 207:34]
  wire  sum_3902 = sum_3829 ^ cout_3828; // @[Mul.scala 206:34]
  wire  sum_3947 = sum_3874 ^ cout_3873; // @[Mul.scala 206:34]
  wire  cout_3947 = sum_3874 & cout_3873; // @[Mul.scala 207:34]
  wire  sum_3948 = sum_3875 ^ cout_3874; // @[Mul.scala 206:34]
  wire  cout_3948 = sum_3875 & cout_3874; // @[Mul.scala 207:34]
  wire  sum_3949 = sum_3876 ^ cout_3875; // @[Mul.scala 206:34]
  wire  cout_3949 = sum_3876 & cout_3875; // @[Mul.scala 207:34]
  wire  _sum_T_4635 = sum_3877 ^ sum_3878; // @[Mul.scala 191:34]
  wire  sum_3950 = sum_3877 ^ sum_3878 ^ cout_3876; // @[Mul.scala 191:42]
  wire  cout_3950 = sum_3877 & sum_3878 | _sum_T_4635 & cout_3876; // @[Mul.scala 192:44]
  wire  sum_3951 = sum_3879 ^ sum_3880; // @[Mul.scala 206:34]
  wire  cout_3951 = sum_3879 & sum_3880; // @[Mul.scala 207:34]
  wire  sum_3952 = cout_3877 ^ cout_3878; // @[Mul.scala 206:34]
  wire  cout_3952 = cout_3877 & cout_3878; // @[Mul.scala 207:34]
  wire  sum_3953 = sum_3881 ^ sum_3882; // @[Mul.scala 206:34]
  wire  cout_3953 = sum_3881 & sum_3882; // @[Mul.scala 207:34]
  wire  sum_3954 = cout_3879 ^ cout_3880; // @[Mul.scala 206:34]
  wire  cout_3954 = cout_3879 & cout_3880; // @[Mul.scala 207:34]
  wire  sum_3955 = sum_3883 ^ sum_3884; // @[Mul.scala 206:34]
  wire  cout_3955 = sum_3883 & sum_3884; // @[Mul.scala 207:34]
  wire  sum_3956 = cout_3881 ^ cout_3882; // @[Mul.scala 206:34]
  wire  cout_3956 = cout_3881 & cout_3882; // @[Mul.scala 207:34]
  wire  sum_3957 = sum_3885 ^ sum_3886; // @[Mul.scala 206:34]
  wire  cout_3957 = sum_3885 & sum_3886; // @[Mul.scala 207:34]
  wire  sum_3958 = cout_3883 ^ cout_3884; // @[Mul.scala 206:34]
  wire  cout_3958 = cout_3883 & cout_3884; // @[Mul.scala 207:34]
  wire  sum_3959 = sum_3887 ^ sum_3888; // @[Mul.scala 206:34]
  wire  cout_3959 = sum_3887 & sum_3888; // @[Mul.scala 207:34]
  wire  sum_3960 = cout_3885 ^ cout_3886; // @[Mul.scala 206:34]
  wire  cout_3960 = cout_3885 & cout_3886; // @[Mul.scala 207:34]
  wire  sum_3961 = sum_3889 ^ sum_3890; // @[Mul.scala 206:34]
  wire  cout_3961 = sum_3889 & sum_3890; // @[Mul.scala 207:34]
  wire  sum_3962 = cout_3887 ^ cout_3888; // @[Mul.scala 206:34]
  wire  cout_3962 = cout_3887 & cout_3888; // @[Mul.scala 207:34]
  wire  sum_3963 = sum_3891 ^ sum_3892; // @[Mul.scala 206:34]
  wire  cout_3963 = sum_3891 & sum_3892; // @[Mul.scala 207:34]
  wire  sum_3964 = cout_3889 ^ cout_3890; // @[Mul.scala 206:34]
  wire  cout_3964 = cout_3889 & cout_3890; // @[Mul.scala 207:34]
  wire  sum_3965 = sum_3893 ^ sum_3894; // @[Mul.scala 206:34]
  wire  cout_3965 = sum_3893 & sum_3894; // @[Mul.scala 207:34]
  wire  sum_3966 = cout_3891 ^ cout_3892; // @[Mul.scala 206:34]
  wire  cout_3966 = cout_3891 & cout_3892; // @[Mul.scala 207:34]
  wire  sum_3967 = sum_3895 ^ sum_3896; // @[Mul.scala 206:34]
  wire  cout_3967 = sum_3895 & sum_3896; // @[Mul.scala 207:34]
  wire  sum_3968 = cout_3893 ^ cout_3894; // @[Mul.scala 206:34]
  wire  cout_3968 = cout_3893 & cout_3894; // @[Mul.scala 207:34]
  wire  _sum_T_4655 = sum_3897 ^ cout_3895; // @[Mul.scala 191:34]
  wire  sum_3969 = sum_3897 ^ cout_3895 ^ cout_3896; // @[Mul.scala 191:42]
  wire  cout_3969 = sum_3897 & cout_3895 | _sum_T_4655 & cout_3896; // @[Mul.scala 192:44]
  wire  sum_3970 = sum_3898 ^ cout_3897; // @[Mul.scala 206:34]
  wire  cout_3970 = sum_3898 & cout_3897; // @[Mul.scala 207:34]
  wire  sum_3971 = sum_3899 ^ cout_3898; // @[Mul.scala 206:34]
  wire  cout_3971 = sum_3899 & cout_3898; // @[Mul.scala 207:34]
  wire  sum_3972 = sum_3900 ^ cout_3899; // @[Mul.scala 206:34]
  wire  cout_3972 = sum_3900 & cout_3899; // @[Mul.scala 207:34]
  wire  sum_3973 = sum_3901 ^ cout_3900; // @[Mul.scala 206:34]
  wire  cout_3973 = sum_3901 & cout_3900; // @[Mul.scala 207:34]
  wire  sum_3974 = sum_3902 ^ cout_3901; // @[Mul.scala 206:34]
  wire  sum_4020 = sum_3948 ^ cout_3947; // @[Mul.scala 206:34]
  wire  cout_4020 = sum_3948 & cout_3947; // @[Mul.scala 207:34]
  wire  sum_4021 = sum_3949 ^ cout_3948; // @[Mul.scala 206:34]
  wire  cout_4021 = sum_3949 & cout_3948; // @[Mul.scala 207:34]
  wire  sum_4022 = sum_3950 ^ cout_3949; // @[Mul.scala 206:34]
  wire  cout_4022 = sum_3950 & cout_3949; // @[Mul.scala 207:34]
  wire  _sum_T_4710 = sum_3951 ^ sum_3952; // @[Mul.scala 191:34]
  wire  sum_4023 = sum_3951 ^ sum_3952 ^ cout_3950; // @[Mul.scala 191:42]
  wire  cout_4023 = sum_3951 & sum_3952 | _sum_T_4710 & cout_3950; // @[Mul.scala 192:44]
  wire  sum_4024 = sum_3953 ^ sum_3954; // @[Mul.scala 206:34]
  wire  cout_4024 = sum_3953 & sum_3954; // @[Mul.scala 207:34]
  wire  sum_4025 = cout_3951 ^ cout_3952; // @[Mul.scala 206:34]
  wire  cout_4025 = cout_3951 & cout_3952; // @[Mul.scala 207:34]
  wire  sum_4026 = sum_3955 ^ sum_3956; // @[Mul.scala 206:34]
  wire  cout_4026 = sum_3955 & sum_3956; // @[Mul.scala 207:34]
  wire  sum_4027 = cout_3953 ^ cout_3954; // @[Mul.scala 206:34]
  wire  cout_4027 = cout_3953 & cout_3954; // @[Mul.scala 207:34]
  wire  sum_4028 = sum_3957 ^ sum_3958; // @[Mul.scala 206:34]
  wire  cout_4028 = sum_3957 & sum_3958; // @[Mul.scala 207:34]
  wire  sum_4029 = cout_3955 ^ cout_3956; // @[Mul.scala 206:34]
  wire  cout_4029 = cout_3955 & cout_3956; // @[Mul.scala 207:34]
  wire  sum_4030 = sum_3959 ^ sum_3960; // @[Mul.scala 206:34]
  wire  cout_4030 = sum_3959 & sum_3960; // @[Mul.scala 207:34]
  wire  sum_4031 = cout_3957 ^ cout_3958; // @[Mul.scala 206:34]
  wire  cout_4031 = cout_3957 & cout_3958; // @[Mul.scala 207:34]
  wire  sum_4032 = sum_3961 ^ sum_3962; // @[Mul.scala 206:34]
  wire  cout_4032 = sum_3961 & sum_3962; // @[Mul.scala 207:34]
  wire  sum_4033 = cout_3959 ^ cout_3960; // @[Mul.scala 206:34]
  wire  cout_4033 = cout_3959 & cout_3960; // @[Mul.scala 207:34]
  wire  sum_4034 = sum_3963 ^ sum_3964; // @[Mul.scala 206:34]
  wire  cout_4034 = sum_3963 & sum_3964; // @[Mul.scala 207:34]
  wire  sum_4035 = cout_3961 ^ cout_3962; // @[Mul.scala 206:34]
  wire  cout_4035 = cout_3961 & cout_3962; // @[Mul.scala 207:34]
  wire  sum_4036 = sum_3965 ^ sum_3966; // @[Mul.scala 206:34]
  wire  cout_4036 = sum_3965 & sum_3966; // @[Mul.scala 207:34]
  wire  sum_4037 = cout_3963 ^ cout_3964; // @[Mul.scala 206:34]
  wire  cout_4037 = cout_3963 & cout_3964; // @[Mul.scala 207:34]
  wire  sum_4038 = sum_3967 ^ sum_3968; // @[Mul.scala 206:34]
  wire  cout_4038 = sum_3967 & sum_3968; // @[Mul.scala 207:34]
  wire  sum_4039 = cout_3965 ^ cout_3966; // @[Mul.scala 206:34]
  wire  cout_4039 = cout_3965 & cout_3966; // @[Mul.scala 207:34]
  wire  _sum_T_4728 = sum_3969 ^ cout_3967; // @[Mul.scala 191:34]
  wire  sum_4040 = sum_3969 ^ cout_3967 ^ cout_3968; // @[Mul.scala 191:42]
  wire  cout_4040 = sum_3969 & cout_3967 | _sum_T_4728 & cout_3968; // @[Mul.scala 192:44]
  wire  sum_4041 = sum_3970 ^ cout_3969; // @[Mul.scala 206:34]
  wire  cout_4041 = sum_3970 & cout_3969; // @[Mul.scala 207:34]
  wire  sum_4042 = sum_3971 ^ cout_3970; // @[Mul.scala 206:34]
  wire  cout_4042 = sum_3971 & cout_3970; // @[Mul.scala 207:34]
  wire  sum_4043 = sum_3972 ^ cout_3971; // @[Mul.scala 206:34]
  wire  cout_4043 = sum_3972 & cout_3971; // @[Mul.scala 207:34]
  wire  sum_4044 = sum_3973 ^ cout_3972; // @[Mul.scala 206:34]
  wire  cout_4044 = sum_3973 & cout_3972; // @[Mul.scala 207:34]
  wire  sum_4045 = sum_3974 ^ cout_3973; // @[Mul.scala 206:34]
  wire  sum_4092 = sum_4021 ^ cout_4020; // @[Mul.scala 206:34]
  wire  cout_4092 = sum_4021 & cout_4020; // @[Mul.scala 207:34]
  wire  sum_4093 = sum_4022 ^ cout_4021; // @[Mul.scala 206:34]
  wire  cout_4093 = sum_4022 & cout_4021; // @[Mul.scala 207:34]
  wire  sum_4094 = sum_4023 ^ cout_4022; // @[Mul.scala 206:34]
  wire  cout_4094 = sum_4023 & cout_4022; // @[Mul.scala 207:34]
  wire  _sum_T_4784 = sum_4024 ^ sum_4025; // @[Mul.scala 191:34]
  wire  sum_4095 = sum_4024 ^ sum_4025 ^ cout_4023; // @[Mul.scala 191:42]
  wire  cout_4095 = sum_4024 & sum_4025 | _sum_T_4784 & cout_4023; // @[Mul.scala 192:44]
  wire  sum_4096 = sum_4026 ^ sum_4027; // @[Mul.scala 206:34]
  wire  cout_4096 = sum_4026 & sum_4027; // @[Mul.scala 207:34]
  wire  sum_4097 = cout_4024 ^ cout_4025; // @[Mul.scala 206:34]
  wire  cout_4097 = cout_4024 & cout_4025; // @[Mul.scala 207:34]
  wire  sum_4098 = sum_4028 ^ sum_4029; // @[Mul.scala 206:34]
  wire  cout_4098 = sum_4028 & sum_4029; // @[Mul.scala 207:34]
  wire  sum_4099 = cout_4026 ^ cout_4027; // @[Mul.scala 206:34]
  wire  cout_4099 = cout_4026 & cout_4027; // @[Mul.scala 207:34]
  wire  sum_4100 = sum_4030 ^ sum_4031; // @[Mul.scala 206:34]
  wire  cout_4100 = sum_4030 & sum_4031; // @[Mul.scala 207:34]
  wire  sum_4101 = cout_4028 ^ cout_4029; // @[Mul.scala 206:34]
  wire  cout_4101 = cout_4028 & cout_4029; // @[Mul.scala 207:34]
  wire  sum_4102 = sum_4032 ^ sum_4033; // @[Mul.scala 206:34]
  wire  cout_4102 = sum_4032 & sum_4033; // @[Mul.scala 207:34]
  wire  sum_4103 = cout_4030 ^ cout_4031; // @[Mul.scala 206:34]
  wire  cout_4103 = cout_4030 & cout_4031; // @[Mul.scala 207:34]
  wire  sum_4104 = sum_4034 ^ sum_4035; // @[Mul.scala 206:34]
  wire  cout_4104 = sum_4034 & sum_4035; // @[Mul.scala 207:34]
  wire  sum_4105 = cout_4032 ^ cout_4033; // @[Mul.scala 206:34]
  wire  cout_4105 = cout_4032 & cout_4033; // @[Mul.scala 207:34]
  wire  sum_4106 = sum_4036 ^ sum_4037; // @[Mul.scala 206:34]
  wire  cout_4106 = sum_4036 & sum_4037; // @[Mul.scala 207:34]
  wire  sum_4107 = cout_4034 ^ cout_4035; // @[Mul.scala 206:34]
  wire  cout_4107 = cout_4034 & cout_4035; // @[Mul.scala 207:34]
  wire  sum_4108 = sum_4038 ^ sum_4039; // @[Mul.scala 206:34]
  wire  cout_4108 = sum_4038 & sum_4039; // @[Mul.scala 207:34]
  wire  sum_4109 = cout_4036 ^ cout_4037; // @[Mul.scala 206:34]
  wire  cout_4109 = cout_4036 & cout_4037; // @[Mul.scala 207:34]
  wire  _sum_T_4800 = sum_4040 ^ cout_4038; // @[Mul.scala 191:34]
  wire  sum_4110 = sum_4040 ^ cout_4038 ^ cout_4039; // @[Mul.scala 191:42]
  wire  cout_4110 = sum_4040 & cout_4038 | _sum_T_4800 & cout_4039; // @[Mul.scala 192:44]
  wire  sum_4111 = sum_4041 ^ cout_4040; // @[Mul.scala 206:34]
  wire  cout_4111 = sum_4041 & cout_4040; // @[Mul.scala 207:34]
  wire  sum_4112 = sum_4042 ^ cout_4041; // @[Mul.scala 206:34]
  wire  cout_4112 = sum_4042 & cout_4041; // @[Mul.scala 207:34]
  wire  sum_4113 = sum_4043 ^ cout_4042; // @[Mul.scala 206:34]
  wire  cout_4113 = sum_4043 & cout_4042; // @[Mul.scala 207:34]
  wire  sum_4114 = sum_4044 ^ cout_4043; // @[Mul.scala 206:34]
  wire  cout_4114 = sum_4044 & cout_4043; // @[Mul.scala 207:34]
  wire  sum_4115 = sum_4045 ^ cout_4044; // @[Mul.scala 206:34]
  wire  sum_4163 = sum_4093 ^ cout_4092; // @[Mul.scala 206:34]
  wire  cout_4163 = sum_4093 & cout_4092; // @[Mul.scala 207:34]
  wire  sum_4164 = sum_4094 ^ cout_4093; // @[Mul.scala 206:34]
  wire  cout_4164 = sum_4094 & cout_4093; // @[Mul.scala 207:34]
  wire  sum_4165 = sum_4095 ^ cout_4094; // @[Mul.scala 206:34]
  wire  cout_4165 = sum_4095 & cout_4094; // @[Mul.scala 207:34]
  wire  _sum_T_4857 = sum_4096 ^ sum_4097; // @[Mul.scala 191:34]
  wire  sum_4166 = sum_4096 ^ sum_4097 ^ cout_4095; // @[Mul.scala 191:42]
  wire  cout_4166 = sum_4096 & sum_4097 | _sum_T_4857 & cout_4095; // @[Mul.scala 192:44]
  wire  sum_4167 = sum_4098 ^ sum_4099; // @[Mul.scala 206:34]
  wire  cout_4167 = sum_4098 & sum_4099; // @[Mul.scala 207:34]
  wire  sum_4168 = cout_4096 ^ cout_4097; // @[Mul.scala 206:34]
  wire  cout_4168 = cout_4096 & cout_4097; // @[Mul.scala 207:34]
  wire  sum_4169 = sum_4100 ^ sum_4101; // @[Mul.scala 206:34]
  wire  cout_4169 = sum_4100 & sum_4101; // @[Mul.scala 207:34]
  wire  sum_4170 = cout_4098 ^ cout_4099; // @[Mul.scala 206:34]
  wire  cout_4170 = cout_4098 & cout_4099; // @[Mul.scala 207:34]
  wire  sum_4171 = sum_4102 ^ sum_4103; // @[Mul.scala 206:34]
  wire  cout_4171 = sum_4102 & sum_4103; // @[Mul.scala 207:34]
  wire  sum_4172 = cout_4100 ^ cout_4101; // @[Mul.scala 206:34]
  wire  cout_4172 = cout_4100 & cout_4101; // @[Mul.scala 207:34]
  wire  sum_4173 = sum_4104 ^ sum_4105; // @[Mul.scala 206:34]
  wire  cout_4173 = sum_4104 & sum_4105; // @[Mul.scala 207:34]
  wire  sum_4174 = cout_4102 ^ cout_4103; // @[Mul.scala 206:34]
  wire  cout_4174 = cout_4102 & cout_4103; // @[Mul.scala 207:34]
  wire  sum_4175 = sum_4106 ^ sum_4107; // @[Mul.scala 206:34]
  wire  cout_4175 = sum_4106 & sum_4107; // @[Mul.scala 207:34]
  wire  sum_4176 = cout_4104 ^ cout_4105; // @[Mul.scala 206:34]
  wire  cout_4176 = cout_4104 & cout_4105; // @[Mul.scala 207:34]
  wire  sum_4177 = sum_4108 ^ sum_4109; // @[Mul.scala 206:34]
  wire  cout_4177 = sum_4108 & sum_4109; // @[Mul.scala 207:34]
  wire  sum_4178 = cout_4106 ^ cout_4107; // @[Mul.scala 206:34]
  wire  cout_4178 = cout_4106 & cout_4107; // @[Mul.scala 207:34]
  wire  _sum_T_4871 = sum_4110 ^ cout_4108; // @[Mul.scala 191:34]
  wire  sum_4179 = sum_4110 ^ cout_4108 ^ cout_4109; // @[Mul.scala 191:42]
  wire  cout_4179 = sum_4110 & cout_4108 | _sum_T_4871 & cout_4109; // @[Mul.scala 192:44]
  wire  sum_4180 = sum_4111 ^ cout_4110; // @[Mul.scala 206:34]
  wire  cout_4180 = sum_4111 & cout_4110; // @[Mul.scala 207:34]
  wire  sum_4181 = sum_4112 ^ cout_4111; // @[Mul.scala 206:34]
  wire  cout_4181 = sum_4112 & cout_4111; // @[Mul.scala 207:34]
  wire  sum_4182 = sum_4113 ^ cout_4112; // @[Mul.scala 206:34]
  wire  cout_4182 = sum_4113 & cout_4112; // @[Mul.scala 207:34]
  wire  sum_4183 = sum_4114 ^ cout_4113; // @[Mul.scala 206:34]
  wire  cout_4183 = sum_4114 & cout_4113; // @[Mul.scala 207:34]
  wire  sum_4184 = sum_4115 ^ cout_4114; // @[Mul.scala 206:34]
  wire  sum_4233 = sum_4164 ^ cout_4163; // @[Mul.scala 206:34]
  wire  cout_4233 = sum_4164 & cout_4163; // @[Mul.scala 207:34]
  wire  sum_4234 = sum_4165 ^ cout_4164; // @[Mul.scala 206:34]
  wire  cout_4234 = sum_4165 & cout_4164; // @[Mul.scala 207:34]
  wire  sum_4235 = sum_4166 ^ cout_4165; // @[Mul.scala 206:34]
  wire  cout_4235 = sum_4166 & cout_4165; // @[Mul.scala 207:34]
  wire  _sum_T_4929 = sum_4167 ^ sum_4168; // @[Mul.scala 191:34]
  wire  sum_4236 = sum_4167 ^ sum_4168 ^ cout_4166; // @[Mul.scala 191:42]
  wire  cout_4236 = sum_4167 & sum_4168 | _sum_T_4929 & cout_4166; // @[Mul.scala 192:44]
  wire  sum_4237 = sum_4169 ^ sum_4170; // @[Mul.scala 206:34]
  wire  cout_4237 = sum_4169 & sum_4170; // @[Mul.scala 207:34]
  wire  sum_4238 = cout_4167 ^ cout_4168; // @[Mul.scala 206:34]
  wire  cout_4238 = cout_4167 & cout_4168; // @[Mul.scala 207:34]
  wire  sum_4239 = sum_4171 ^ sum_4172; // @[Mul.scala 206:34]
  wire  cout_4239 = sum_4171 & sum_4172; // @[Mul.scala 207:34]
  wire  sum_4240 = cout_4169 ^ cout_4170; // @[Mul.scala 206:34]
  wire  cout_4240 = cout_4169 & cout_4170; // @[Mul.scala 207:34]
  wire  sum_4241 = sum_4173 ^ sum_4174; // @[Mul.scala 206:34]
  wire  cout_4241 = sum_4173 & sum_4174; // @[Mul.scala 207:34]
  wire  sum_4242 = cout_4171 ^ cout_4172; // @[Mul.scala 206:34]
  wire  cout_4242 = cout_4171 & cout_4172; // @[Mul.scala 207:34]
  wire  sum_4243 = sum_4175 ^ sum_4176; // @[Mul.scala 206:34]
  wire  cout_4243 = sum_4175 & sum_4176; // @[Mul.scala 207:34]
  wire  sum_4244 = cout_4173 ^ cout_4174; // @[Mul.scala 206:34]
  wire  cout_4244 = cout_4173 & cout_4174; // @[Mul.scala 207:34]
  wire  sum_4245 = sum_4177 ^ sum_4178; // @[Mul.scala 206:34]
  wire  cout_4245 = sum_4177 & sum_4178; // @[Mul.scala 207:34]
  wire  sum_4246 = cout_4175 ^ cout_4176; // @[Mul.scala 206:34]
  wire  cout_4246 = cout_4175 & cout_4176; // @[Mul.scala 207:34]
  wire  _sum_T_4941 = sum_4179 ^ cout_4177; // @[Mul.scala 191:34]
  wire  sum_4247 = sum_4179 ^ cout_4177 ^ cout_4178; // @[Mul.scala 191:42]
  wire  cout_4247 = sum_4179 & cout_4177 | _sum_T_4941 & cout_4178; // @[Mul.scala 192:44]
  wire  sum_4248 = sum_4180 ^ cout_4179; // @[Mul.scala 206:34]
  wire  cout_4248 = sum_4180 & cout_4179; // @[Mul.scala 207:34]
  wire  sum_4249 = sum_4181 ^ cout_4180; // @[Mul.scala 206:34]
  wire  cout_4249 = sum_4181 & cout_4180; // @[Mul.scala 207:34]
  wire  sum_4250 = sum_4182 ^ cout_4181; // @[Mul.scala 206:34]
  wire  cout_4250 = sum_4182 & cout_4181; // @[Mul.scala 207:34]
  wire  sum_4251 = sum_4183 ^ cout_4182; // @[Mul.scala 206:34]
  wire  cout_4251 = sum_4183 & cout_4182; // @[Mul.scala 207:34]
  wire  sum_4252 = sum_4184 ^ cout_4183; // @[Mul.scala 206:34]
  wire  sum_4302 = sum_4234 ^ cout_4233; // @[Mul.scala 206:34]
  wire  cout_4302 = sum_4234 & cout_4233; // @[Mul.scala 207:34]
  wire  sum_4303 = sum_4235 ^ cout_4234; // @[Mul.scala 206:34]
  wire  cout_4303 = sum_4235 & cout_4234; // @[Mul.scala 207:34]
  wire  sum_4304 = sum_4236 ^ cout_4235; // @[Mul.scala 206:34]
  wire  cout_4304 = sum_4236 & cout_4235; // @[Mul.scala 207:34]
  wire  _sum_T_5000 = sum_4237 ^ sum_4238; // @[Mul.scala 191:34]
  wire  sum_4305 = sum_4237 ^ sum_4238 ^ cout_4236; // @[Mul.scala 191:42]
  wire  cout_4305 = sum_4237 & sum_4238 | _sum_T_5000 & cout_4236; // @[Mul.scala 192:44]
  wire  sum_4306 = sum_4239 ^ sum_4240; // @[Mul.scala 206:34]
  wire  cout_4306 = sum_4239 & sum_4240; // @[Mul.scala 207:34]
  wire  sum_4307 = cout_4237 ^ cout_4238; // @[Mul.scala 206:34]
  wire  cout_4307 = cout_4237 & cout_4238; // @[Mul.scala 207:34]
  wire  sum_4308 = sum_4241 ^ sum_4242; // @[Mul.scala 206:34]
  wire  cout_4308 = sum_4241 & sum_4242; // @[Mul.scala 207:34]
  wire  sum_4309 = cout_4239 ^ cout_4240; // @[Mul.scala 206:34]
  wire  cout_4309 = cout_4239 & cout_4240; // @[Mul.scala 207:34]
  wire  sum_4310 = sum_4243 ^ sum_4244; // @[Mul.scala 206:34]
  wire  cout_4310 = sum_4243 & sum_4244; // @[Mul.scala 207:34]
  wire  sum_4311 = cout_4241 ^ cout_4242; // @[Mul.scala 206:34]
  wire  cout_4311 = cout_4241 & cout_4242; // @[Mul.scala 207:34]
  wire  sum_4312 = sum_4245 ^ sum_4246; // @[Mul.scala 206:34]
  wire  cout_4312 = sum_4245 & sum_4246; // @[Mul.scala 207:34]
  wire  sum_4313 = cout_4243 ^ cout_4244; // @[Mul.scala 206:34]
  wire  cout_4313 = cout_4243 & cout_4244; // @[Mul.scala 207:34]
  wire  _sum_T_5010 = sum_4247 ^ cout_4245; // @[Mul.scala 191:34]
  wire  sum_4314 = sum_4247 ^ cout_4245 ^ cout_4246; // @[Mul.scala 191:42]
  wire  cout_4314 = sum_4247 & cout_4245 | _sum_T_5010 & cout_4246; // @[Mul.scala 192:44]
  wire  sum_4315 = sum_4248 ^ cout_4247; // @[Mul.scala 206:34]
  wire  cout_4315 = sum_4248 & cout_4247; // @[Mul.scala 207:34]
  wire  sum_4316 = sum_4249 ^ cout_4248; // @[Mul.scala 206:34]
  wire  cout_4316 = sum_4249 & cout_4248; // @[Mul.scala 207:34]
  wire  sum_4317 = sum_4250 ^ cout_4249; // @[Mul.scala 206:34]
  wire  cout_4317 = sum_4250 & cout_4249; // @[Mul.scala 207:34]
  wire  sum_4318 = sum_4251 ^ cout_4250; // @[Mul.scala 206:34]
  wire  cout_4318 = sum_4251 & cout_4250; // @[Mul.scala 207:34]
  wire  sum_4319 = sum_4252 ^ cout_4251; // @[Mul.scala 206:34]
  wire  sum_4370 = sum_4303 ^ cout_4302; // @[Mul.scala 206:34]
  wire  cout_4370 = sum_4303 & cout_4302; // @[Mul.scala 207:34]
  wire  sum_4371 = sum_4304 ^ cout_4303; // @[Mul.scala 206:34]
  wire  cout_4371 = sum_4304 & cout_4303; // @[Mul.scala 207:34]
  wire  sum_4372 = sum_4305 ^ cout_4304; // @[Mul.scala 206:34]
  wire  cout_4372 = sum_4305 & cout_4304; // @[Mul.scala 207:34]
  wire  _sum_T_5070 = sum_4306 ^ sum_4307; // @[Mul.scala 191:34]
  wire  sum_4373 = sum_4306 ^ sum_4307 ^ cout_4305; // @[Mul.scala 191:42]
  wire  cout_4373 = sum_4306 & sum_4307 | _sum_T_5070 & cout_4305; // @[Mul.scala 192:44]
  wire  sum_4374 = sum_4308 ^ sum_4309; // @[Mul.scala 206:34]
  wire  cout_4374 = sum_4308 & sum_4309; // @[Mul.scala 207:34]
  wire  sum_4375 = cout_4306 ^ cout_4307; // @[Mul.scala 206:34]
  wire  cout_4375 = cout_4306 & cout_4307; // @[Mul.scala 207:34]
  wire  sum_4376 = sum_4310 ^ sum_4311; // @[Mul.scala 206:34]
  wire  cout_4376 = sum_4310 & sum_4311; // @[Mul.scala 207:34]
  wire  sum_4377 = cout_4308 ^ cout_4309; // @[Mul.scala 206:34]
  wire  cout_4377 = cout_4308 & cout_4309; // @[Mul.scala 207:34]
  wire  sum_4378 = sum_4312 ^ sum_4313; // @[Mul.scala 206:34]
  wire  cout_4378 = sum_4312 & sum_4313; // @[Mul.scala 207:34]
  wire  sum_4379 = cout_4310 ^ cout_4311; // @[Mul.scala 206:34]
  wire  cout_4379 = cout_4310 & cout_4311; // @[Mul.scala 207:34]
  wire  _sum_T_5078 = sum_4314 ^ cout_4312; // @[Mul.scala 191:34]
  wire  sum_4380 = sum_4314 ^ cout_4312 ^ cout_4313; // @[Mul.scala 191:42]
  wire  cout_4380 = sum_4314 & cout_4312 | _sum_T_5078 & cout_4313; // @[Mul.scala 192:44]
  wire  sum_4381 = sum_4315 ^ cout_4314; // @[Mul.scala 206:34]
  wire  cout_4381 = sum_4315 & cout_4314; // @[Mul.scala 207:34]
  wire  sum_4382 = sum_4316 ^ cout_4315; // @[Mul.scala 206:34]
  wire  cout_4382 = sum_4316 & cout_4315; // @[Mul.scala 207:34]
  wire  sum_4383 = sum_4317 ^ cout_4316; // @[Mul.scala 206:34]
  wire  cout_4383 = sum_4317 & cout_4316; // @[Mul.scala 207:34]
  wire  sum_4384 = sum_4318 ^ cout_4317; // @[Mul.scala 206:34]
  wire  cout_4384 = sum_4318 & cout_4317; // @[Mul.scala 207:34]
  wire  sum_4385 = sum_4319 ^ cout_4318; // @[Mul.scala 206:34]
  wire  sum_4437 = sum_4371 ^ cout_4370; // @[Mul.scala 206:34]
  wire  cout_4437 = sum_4371 & cout_4370; // @[Mul.scala 207:34]
  wire  sum_4438 = sum_4372 ^ cout_4371; // @[Mul.scala 206:34]
  wire  cout_4438 = sum_4372 & cout_4371; // @[Mul.scala 207:34]
  wire  sum_4439 = sum_4373 ^ cout_4372; // @[Mul.scala 206:34]
  wire  cout_4439 = sum_4373 & cout_4372; // @[Mul.scala 207:34]
  wire  _sum_T_5139 = sum_4374 ^ sum_4375; // @[Mul.scala 191:34]
  wire  sum_4440 = sum_4374 ^ sum_4375 ^ cout_4373; // @[Mul.scala 191:42]
  wire  cout_4440 = sum_4374 & sum_4375 | _sum_T_5139 & cout_4373; // @[Mul.scala 192:44]
  wire  sum_4441 = sum_4376 ^ sum_4377; // @[Mul.scala 206:34]
  wire  cout_4441 = sum_4376 & sum_4377; // @[Mul.scala 207:34]
  wire  sum_4442 = cout_4374 ^ cout_4375; // @[Mul.scala 206:34]
  wire  cout_4442 = cout_4374 & cout_4375; // @[Mul.scala 207:34]
  wire  sum_4443 = sum_4378 ^ sum_4379; // @[Mul.scala 206:34]
  wire  cout_4443 = sum_4378 & sum_4379; // @[Mul.scala 207:34]
  wire  sum_4444 = cout_4376 ^ cout_4377; // @[Mul.scala 206:34]
  wire  cout_4444 = cout_4376 & cout_4377; // @[Mul.scala 207:34]
  wire  _sum_T_5145 = sum_4380 ^ cout_4378; // @[Mul.scala 191:34]
  wire  sum_4445 = sum_4380 ^ cout_4378 ^ cout_4379; // @[Mul.scala 191:42]
  wire  cout_4445 = sum_4380 & cout_4378 | _sum_T_5145 & cout_4379; // @[Mul.scala 192:44]
  wire  sum_4446 = sum_4381 ^ cout_4380; // @[Mul.scala 206:34]
  wire  cout_4446 = sum_4381 & cout_4380; // @[Mul.scala 207:34]
  wire  sum_4447 = sum_4382 ^ cout_4381; // @[Mul.scala 206:34]
  wire  cout_4447 = sum_4382 & cout_4381; // @[Mul.scala 207:34]
  wire  sum_4448 = sum_4383 ^ cout_4382; // @[Mul.scala 206:34]
  wire  cout_4448 = sum_4383 & cout_4382; // @[Mul.scala 207:34]
  wire  sum_4449 = sum_4384 ^ cout_4383; // @[Mul.scala 206:34]
  wire  cout_4449 = sum_4384 & cout_4383; // @[Mul.scala 207:34]
  wire  sum_4450 = sum_4385 ^ cout_4384; // @[Mul.scala 206:34]
  wire  sum_4503 = sum_4438 ^ cout_4437; // @[Mul.scala 206:34]
  wire  cout_4503 = sum_4438 & cout_4437; // @[Mul.scala 207:34]
  wire  sum_4504 = sum_4439 ^ cout_4438; // @[Mul.scala 206:34]
  wire  cout_4504 = sum_4439 & cout_4438; // @[Mul.scala 207:34]
  wire  sum_4505 = sum_4440 ^ cout_4439; // @[Mul.scala 206:34]
  wire  cout_4505 = sum_4440 & cout_4439; // @[Mul.scala 207:34]
  wire  _sum_T_5207 = sum_4441 ^ sum_4442; // @[Mul.scala 191:34]
  wire  sum_4506 = sum_4441 ^ sum_4442 ^ cout_4440; // @[Mul.scala 191:42]
  wire  cout_4506 = sum_4441 & sum_4442 | _sum_T_5207 & cout_4440; // @[Mul.scala 192:44]
  wire  sum_4507 = sum_4443 ^ sum_4444; // @[Mul.scala 206:34]
  wire  cout_4507 = sum_4443 & sum_4444; // @[Mul.scala 207:34]
  wire  sum_4508 = cout_4441 ^ cout_4442; // @[Mul.scala 206:34]
  wire  cout_4508 = cout_4441 & cout_4442; // @[Mul.scala 207:34]
  wire  _sum_T_5211 = sum_4445 ^ cout_4443; // @[Mul.scala 191:34]
  wire  sum_4509 = sum_4445 ^ cout_4443 ^ cout_4444; // @[Mul.scala 191:42]
  wire  cout_4509 = sum_4445 & cout_4443 | _sum_T_5211 & cout_4444; // @[Mul.scala 192:44]
  wire  sum_4510 = sum_4446 ^ cout_4445; // @[Mul.scala 206:34]
  wire  cout_4510 = sum_4446 & cout_4445; // @[Mul.scala 207:34]
  wire  sum_4511 = sum_4447 ^ cout_4446; // @[Mul.scala 206:34]
  wire  cout_4511 = sum_4447 & cout_4446; // @[Mul.scala 207:34]
  wire  sum_4512 = sum_4448 ^ cout_4447; // @[Mul.scala 206:34]
  wire  cout_4512 = sum_4448 & cout_4447; // @[Mul.scala 207:34]
  wire  sum_4513 = sum_4449 ^ cout_4448; // @[Mul.scala 206:34]
  wire  cout_4513 = sum_4449 & cout_4448; // @[Mul.scala 207:34]
  wire  sum_4514 = sum_4450 ^ cout_4449; // @[Mul.scala 206:34]
  wire  sum_4568 = sum_4504 ^ cout_4503; // @[Mul.scala 206:34]
  wire  cout_4568 = sum_4504 & cout_4503; // @[Mul.scala 207:34]
  wire  sum_4569 = sum_4505 ^ cout_4504; // @[Mul.scala 206:34]
  wire  cout_4569 = sum_4505 & cout_4504; // @[Mul.scala 207:34]
  wire  sum_4570 = sum_4506 ^ cout_4505; // @[Mul.scala 206:34]
  wire  cout_4570 = sum_4506 & cout_4505; // @[Mul.scala 207:34]
  wire  _sum_T_5274 = sum_4507 ^ sum_4508; // @[Mul.scala 191:34]
  wire  sum_4571 = sum_4507 ^ sum_4508 ^ cout_4506; // @[Mul.scala 191:42]
  wire  cout_4571 = sum_4507 & sum_4508 | _sum_T_5274 & cout_4506; // @[Mul.scala 192:44]
  wire  _sum_T_5276 = sum_4509 ^ cout_4507; // @[Mul.scala 191:34]
  wire  sum_4572 = sum_4509 ^ cout_4507 ^ cout_4508; // @[Mul.scala 191:42]
  wire  cout_4572 = sum_4509 & cout_4507 | _sum_T_5276 & cout_4508; // @[Mul.scala 192:44]
  wire  sum_4573 = sum_4510 ^ cout_4509; // @[Mul.scala 206:34]
  wire  cout_4573 = sum_4510 & cout_4509; // @[Mul.scala 207:34]
  wire  sum_4574 = sum_4511 ^ cout_4510; // @[Mul.scala 206:34]
  wire  cout_4574 = sum_4511 & cout_4510; // @[Mul.scala 207:34]
  wire  sum_4575 = sum_4512 ^ cout_4511; // @[Mul.scala 206:34]
  wire  cout_4575 = sum_4512 & cout_4511; // @[Mul.scala 207:34]
  wire  sum_4576 = sum_4513 ^ cout_4512; // @[Mul.scala 206:34]
  wire  cout_4576 = sum_4513 & cout_4512; // @[Mul.scala 207:34]
  wire  sum_4577 = sum_4514 ^ cout_4513; // @[Mul.scala 206:34]
  wire [7:0] hi_hi_lo = {cout_4568,1'h0,2'h0,4'h0}; // @[Mul.scala 285:38]
  wire [31:0] hi = {cout_4576,cout_4575,cout_4574,cout_4573,cout_4572,cout_4571,cout_4570,cout_4569,hi_hi_lo,16'h0}; // @[Mul.scala 285:38]
  wire [63:0] _T = {hi,32'h0}; // @[Mul.scala 285:38]
  wire [7:0] lo_lo_lo_1 = {sum_432,sum_320,sum_224,sum_140,sum_66,sum,tree_1_0,tree_0_0}; // @[Mul.scala 285:50]
  wire [15:0] lo_lo_1 = {sum_1292,sum_1188,sum_1083,sum_977,sum_870,sum_762,sum_653,sum_543,lo_lo_lo_1}; // @[Mul.scala 285:50]
  wire [7:0] lo_hi_lo_1 = {sum_2088,sum_1992,sum_1895,sum_1797,sum_1698,sum_1598,sum_1497,sum_1395}; // @[Mul.scala 285:50]
  wire [31:0] lo_1 = {sum_2820,sum_2732,sum_2643,sum_2553,sum_2462,sum_2370,sum_2277,sum_2183,lo_hi_lo_1,lo_lo_1}; // @[Mul.scala 285:50]
  wire [7:0] hi_lo_lo_1 = {sum_3488,sum_3408,sum_3327,sum_3245,sum_3162,sum_3078,sum_2993,sum_2907}; // @[Mul.scala 285:50]
  wire [15:0] hi_lo_1 = {sum_4092,sum_4020,sum_3947,sum_3873,sum_3798,sum_3722,sum_3645,sum_3567,hi_lo_lo_1}; // @[Mul.scala 285:50]
  wire [7:0] hi_hi_lo_1 = {sum_4569,sum_4568,sum_4503,sum_4437,sum_4370,sum_4302,sum_4233,sum_4163}; // @[Mul.scala 285:50]
  wire [31:0] hi_1 = {sum_4577,sum_4576,sum_4575,sum_4574,sum_4573,sum_4572,sum_4571,sum_4570,hi_hi_lo_1,hi_lo_1}; // @[Mul.scala 285:50]
  wire [63:0] _T_1 = {hi_1,lo_1}; // @[Mul.scala 285:50]
  wire  _T_2 = pipeFnlStageInfo_io_enq_ready & pipeFnlStageInfo_io_enq_valid; // @[Decoupled.scala 50:35]
  reg [63:0] sum_4579_0; // @[Reg.scala 16:16]
  reg [63:0] sum_4579_1; // @[Reg.scala 16:16]
  Queue pipeMidStageInfo ( // @[Mul.scala 150:32]
    .clock(pipeMidStageInfo_clock),
    .reset(pipeMidStageInfo_reset),
    .io_enq_ready(pipeMidStageInfo_io_enq_ready),
    .io_enq_valid(pipeMidStageInfo_io_enq_valid),
    .io_enq_bits(pipeMidStageInfo_io_enq_bits),
    .io_deq_ready(pipeMidStageInfo_io_deq_ready),
    .io_deq_valid(pipeMidStageInfo_io_deq_valid),
    .io_deq_bits(pipeMidStageInfo_io_deq_bits)
  );
  Queue pipeFnlStageInfo ( // @[Mul.scala 151:32]
    .clock(pipeFnlStageInfo_clock),
    .reset(pipeFnlStageInfo_reset),
    .io_enq_ready(pipeFnlStageInfo_io_enq_ready),
    .io_enq_valid(pipeFnlStageInfo_io_enq_valid),
    .io_enq_bits(pipeFnlStageInfo_io_enq_bits),
    .io_deq_ready(pipeFnlStageInfo_io_deq_ready),
    .io_deq_valid(pipeFnlStageInfo_io_deq_valid),
    .io_deq_bits(pipeFnlStageInfo_io_deq_bits)
  );
  assign io_enq_ready = pipeMidStageInfo_io_enq_ready; // @[Mul.scala 160:10]
  assign io_deq_valid = pipeFnlStageInfo_io_deq_valid; // @[Mul.scala 162:10]
  assign io_deq_bits = pipeFnlStageInfo_io_deq_bits; // @[Mul.scala 162:10]
  assign io_res = sum_4579_0 + sum_4579_1; // @[Mul.scala 158:21]
  assign pipeMidStageInfo_clock = clock;
  assign pipeMidStageInfo_reset = reset | io_flush; // @[Mul.scala 153:42]
  assign pipeMidStageInfo_io_enq_valid = io_enq_valid; // @[Mul.scala 160:10]
  assign pipeMidStageInfo_io_enq_bits = io_enq_bits; // @[Mul.scala 160:10]
  assign pipeMidStageInfo_io_deq_ready = pipeFnlStageInfo_io_enq_ready; // @[Mul.scala 161:27]
  assign pipeFnlStageInfo_clock = clock;
  assign pipeFnlStageInfo_reset = reset | io_flush; // @[Mul.scala 154:42]
  assign pipeFnlStageInfo_io_enq_valid = pipeMidStageInfo_io_deq_valid; // @[Mul.scala 161:27]
  assign pipeFnlStageInfo_io_enq_bits = pipeMidStageInfo_io_deq_bits; // @[Mul.scala 161:27]
  assign pipeFnlStageInfo_io_deq_ready = io_deq_ready; // @[Mul.scala 162:10]
  always @(posedge clock) begin
    if (_T_2) begin // @[Reg.scala 17:18]
      sum_4579_0 <= _T; // @[Reg.scala 17:22]
    end
    if (_T_2) begin // @[Reg.scala 17:18]
      sum_4579_1 <= _T_1; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  sum_4579_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  sum_4579_1 = _RAND_1[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
